magic
tech sky130A
timestamp 1654536627
<< nwell >>
rect 3509 833 4727 2260
<< nmos >>
rect 3495 505 3895 585
rect 4085 507 4485 587
rect 3495 375 3895 455
rect 4085 377 4485 457
<< pmos >>
rect 3835 1725 4235 2225
rect 3835 1155 4235 1655
rect 4513 1083 4613 1223
rect 3585 898 3785 1068
rect 3835 898 4035 1068
rect 4513 893 4613 1033
<< ndiff >>
rect 3445 573 3495 585
rect 3445 553 3457 573
rect 3477 553 3495 573
rect 3445 505 3495 553
rect 3895 561 3945 585
rect 3895 540 3910 561
rect 3931 540 3945 561
rect 3895 505 3945 540
rect 4035 571 4085 587
rect 4035 550 4051 571
rect 4072 550 4085 571
rect 4035 507 4085 550
rect 4485 561 4535 587
rect 4485 540 4498 561
rect 4519 540 4535 561
rect 4485 507 4535 540
rect 3445 421 3495 455
rect 3445 400 3460 421
rect 3481 400 3495 421
rect 3445 375 3495 400
rect 3895 421 3945 455
rect 3895 400 3910 421
rect 3931 400 3945 421
rect 3895 375 3945 400
rect 4035 421 4085 457
rect 4035 400 4050 421
rect 4071 400 4085 421
rect 4035 377 4085 400
rect 4485 431 4535 457
rect 4485 410 4500 431
rect 4521 410 4535 431
rect 4485 377 4535 410
<< pdiff >>
rect 3785 2198 3835 2225
rect 3785 2177 3800 2198
rect 3821 2177 3835 2198
rect 3785 1725 3835 2177
rect 4235 2203 4285 2225
rect 4235 2182 4248 2203
rect 4269 2182 4285 2203
rect 4235 2050 4285 2182
rect 4235 2000 4257 2050
rect 4278 2000 4285 2050
rect 4235 1766 4285 2000
rect 4235 1745 4249 1766
rect 4270 1745 4285 1766
rect 4235 1725 4285 1745
rect 3785 1206 3835 1655
rect 3785 1185 3800 1206
rect 3821 1185 3835 1206
rect 3785 1155 3835 1185
rect 4235 1641 4285 1655
rect 4235 1620 4249 1641
rect 4270 1620 4285 1641
rect 4235 1155 4285 1620
rect 4463 1143 4513 1223
rect 4463 1122 4476 1143
rect 4497 1122 4513 1143
rect 4463 1083 4513 1122
rect 4613 1214 4663 1223
rect 4613 1193 4627 1214
rect 4648 1193 4663 1214
rect 4613 1110 4663 1193
rect 4613 1089 4626 1110
rect 4647 1089 4663 1110
rect 4613 1083 4663 1089
rect 3535 951 3585 1068
rect 3535 930 3549 951
rect 3570 930 3585 951
rect 3535 898 3585 930
rect 3785 1061 3835 1068
rect 3785 1040 3799 1061
rect 3820 1040 3835 1061
rect 3785 898 3835 1040
rect 4035 941 4085 1068
rect 4035 920 4049 941
rect 4070 920 4085 941
rect 4035 898 4085 920
rect 4463 926 4513 1033
rect 4463 905 4477 926
rect 4498 905 4513 926
rect 4463 893 4513 905
rect 4613 1023 4663 1033
rect 4613 1002 4625 1023
rect 4646 1002 4663 1023
rect 4613 893 4663 1002
<< ndiffc >>
rect 3457 553 3477 573
rect 3910 540 3931 561
rect 4051 550 4072 571
rect 4498 540 4519 561
rect 3460 400 3481 421
rect 3910 400 3931 421
rect 4050 400 4071 421
rect 4500 410 4521 431
<< pdiffc >>
rect 3800 2177 3821 2198
rect 4248 2182 4269 2203
rect 4257 2000 4278 2050
rect 4249 1745 4270 1766
rect 3800 1185 3821 1206
rect 4249 1620 4270 1641
rect 4476 1122 4497 1143
rect 4627 1193 4648 1214
rect 4626 1089 4647 1110
rect 3549 930 3570 951
rect 3799 1040 3820 1061
rect 4049 920 4070 941
rect 4477 905 4498 926
rect 4625 1002 4646 1023
<< psubdiff >>
rect 4535 561 4585 587
rect 4535 539 4544 561
rect 4567 539 4585 561
rect 4535 507 4585 539
<< nsubdiff >>
rect 4285 2050 4335 2225
rect 4285 2000 4295 2050
rect 4316 2000 4335 2050
rect 4285 1725 4335 2000
<< psubdiffcont >>
rect 4544 539 4567 561
<< nsubdiffcont >>
rect 4295 2000 4316 2050
<< poly >>
rect 3870 2295 3940 2310
rect 3870 2265 3890 2295
rect 3920 2265 3940 2295
rect 3870 2255 3940 2265
rect 3835 2225 4235 2255
rect 3835 1655 4235 1725
rect 4524 1292 4565 1298
rect 4524 1271 4533 1292
rect 4554 1271 4565 1292
rect 4524 1248 4565 1271
rect 4513 1223 4613 1248
rect 3835 1135 4235 1155
rect 3585 1068 3785 1093
rect 3835 1068 4035 1093
rect 4513 1033 4613 1083
rect 3585 873 3785 898
rect 3835 873 4035 898
rect 3600 865 3670 873
rect 3600 835 3620 865
rect 3650 835 3670 865
rect 3600 820 3670 835
rect 3850 865 3920 873
rect 4513 868 4613 893
rect 3850 835 3870 865
rect 3900 835 3920 865
rect 3850 820 3920 835
rect 3606 654 3676 668
rect 3606 624 3626 654
rect 3656 624 3676 654
rect 3606 615 3676 624
rect 4120 650 4190 670
rect 4120 620 4140 650
rect 4170 620 4190 650
rect 4120 617 4190 620
rect 3495 585 3895 615
rect 4085 587 4485 617
rect 3495 455 3895 505
rect 4085 457 4485 507
rect 3495 355 3895 375
rect 4085 357 4485 377
<< polycont >>
rect 3890 2265 3920 2295
rect 4533 1271 4554 1292
rect 3620 835 3650 865
rect 3870 835 3900 865
rect 3626 624 3656 654
rect 4140 620 4170 650
<< locali >>
rect 3399 2458 4760 2477
rect 3399 2379 3537 2458
rect 3659 2379 3837 2458
rect 3959 2379 4137 2458
rect 4259 2379 4437 2458
rect 4559 2379 4760 2458
rect 3399 2366 4760 2379
rect 3342 2303 3402 2310
rect 3342 2267 3348 2303
rect 3396 2297 3402 2303
rect 3870 2297 3940 2310
rect 3396 2295 3940 2297
rect 3396 2270 3890 2295
rect 3396 2267 3402 2270
rect 3342 2260 3402 2267
rect 3792 2198 3829 2270
rect 3870 2265 3890 2270
rect 3920 2265 3940 2295
rect 3870 2251 3940 2265
rect 3792 2177 3800 2198
rect 3821 2177 3829 2198
rect 3792 2169 3829 2177
rect 4240 2203 4277 2366
rect 4240 2182 4248 2203
rect 4269 2182 4277 2203
rect 4240 2174 4277 2182
rect 4250 2050 4320 2080
rect 4250 2000 4257 2050
rect 4278 2000 4295 2050
rect 4316 2000 4320 2050
rect 4250 1950 4320 2000
rect 4243 1766 4276 1780
rect 4243 1745 4249 1766
rect 4270 1745 4276 1766
rect 4243 1641 4276 1745
rect 4243 1620 4249 1641
rect 4270 1620 4276 1641
rect 4243 1610 4276 1620
rect 4410 1292 4565 1298
rect 4410 1271 4533 1292
rect 4554 1271 4565 1292
rect 3791 1206 3828 1227
rect 3791 1185 3800 1206
rect 3821 1185 3828 1206
rect 3791 1061 3828 1185
rect 4343 1147 4393 1153
rect 4410 1147 4437 1271
rect 4619 1214 4656 2366
rect 4619 1193 4627 1214
rect 4648 1193 4656 1214
rect 4619 1184 4656 1193
rect 4468 1147 4505 1152
rect 4343 1120 4354 1147
rect 4381 1143 4505 1147
rect 4381 1122 4476 1143
rect 4497 1122 4505 1143
rect 4381 1120 4505 1122
rect 4343 1113 4393 1120
rect 4468 1112 4505 1120
rect 3791 1040 3799 1061
rect 3820 1040 3828 1061
rect 3791 1015 3828 1040
rect 4618 1110 4655 1113
rect 4618 1089 4626 1110
rect 4647 1089 4655 1110
rect 4618 1023 4655 1089
rect 4618 1002 4625 1023
rect 4646 1002 4655 1023
rect 4618 993 4655 1002
rect 3540 954 3580 960
rect 3540 927 3546 954
rect 3573 927 3580 954
rect 3540 920 3580 927
rect 4042 941 4079 960
rect 4042 920 4049 941
rect 4070 920 4079 941
rect 3340 885 3400 892
rect 3340 849 3346 885
rect 3394 881 3400 885
rect 3394 865 3670 881
rect 3394 851 3620 865
rect 3394 849 3400 851
rect 3340 842 3400 849
rect 3600 835 3620 851
rect 3650 835 3670 865
rect 3600 820 3670 835
rect 3850 865 3920 880
rect 3850 835 3870 865
rect 3900 835 3920 865
rect 3850 820 3920 835
rect 3341 801 3401 808
rect 3341 765 3347 801
rect 3395 795 3401 801
rect 3870 795 3900 820
rect 3395 765 3900 795
rect 3341 758 3401 765
rect 3446 736 3489 748
rect 3446 709 3453 736
rect 3480 709 3489 736
rect 3446 700 3489 709
rect 3453 654 3480 700
rect 3606 654 3676 668
rect 3453 624 3626 654
rect 3656 624 3676 654
rect 3453 573 3480 624
rect 3606 608 3676 624
rect 4042 650 4079 920
rect 4470 926 4505 935
rect 4470 905 4477 926
rect 4498 905 4505 926
rect 4470 895 4505 905
rect 4474 860 4501 895
rect 4463 854 4513 860
rect 4463 827 4474 854
rect 4501 827 4513 854
rect 4463 820 4513 827
rect 4120 650 4190 670
rect 4042 620 4140 650
rect 4170 620 4190 650
rect 3453 553 3457 573
rect 3477 553 3480 573
rect 4042 571 4079 620
rect 4120 610 4190 620
rect 3453 530 3480 553
rect 3902 561 3939 570
rect 3902 540 3910 561
rect 3931 540 3939 561
rect 3396 424 3489 430
rect 3396 397 3407 424
rect 3434 421 3489 424
rect 3434 400 3460 421
rect 3481 400 3489 421
rect 3434 397 3489 400
rect 3396 390 3489 397
rect 3902 421 3939 540
rect 4042 550 4051 571
rect 4072 550 4079 571
rect 4042 530 4079 550
rect 4492 561 4573 570
rect 4492 540 4498 561
rect 4519 540 4544 561
rect 4492 539 4544 540
rect 4567 539 4573 561
rect 4492 510 4573 539
rect 4492 431 4529 510
rect 3902 400 3910 421
rect 3931 400 3939 421
rect 3902 286 3939 400
rect 3985 424 4080 430
rect 3985 397 3996 424
rect 4023 421 4080 424
rect 4023 400 4050 421
rect 4071 400 4080 421
rect 4023 397 4080 400
rect 3985 391 4080 397
rect 4492 410 4500 431
rect 4521 410 4529 431
rect 3985 390 4041 391
rect 4492 286 4529 410
rect 3396 268 4759 286
rect 3396 189 3537 268
rect 3659 189 3837 268
rect 3959 189 4137 268
rect 4259 189 4437 268
rect 4559 189 4759 268
rect 3396 177 4759 189
<< viali >>
rect 3537 2379 3659 2458
rect 3837 2379 3959 2458
rect 4137 2379 4259 2458
rect 4437 2379 4559 2458
rect 3348 2267 3396 2303
rect 4354 1120 4381 1147
rect 3546 951 3573 954
rect 3546 930 3549 951
rect 3549 930 3570 951
rect 3570 930 3573 951
rect 3546 927 3573 930
rect 3346 849 3394 885
rect 3347 765 3395 801
rect 3453 709 3480 736
rect 4474 827 4501 854
rect 3407 397 3434 424
rect 3996 397 4023 424
rect 3537 189 3659 268
rect 3837 189 3959 268
rect 4137 189 4259 268
rect 4437 189 4559 268
<< metal1 >>
rect 3399 2458 4760 2477
rect 3399 2379 3537 2458
rect 3659 2379 3837 2458
rect 3959 2379 4137 2458
rect 4259 2379 4437 2458
rect 4559 2379 4760 2458
rect 3399 2366 4760 2379
rect 3342 2303 3402 2310
rect 3342 2267 3348 2303
rect 3396 2267 3402 2303
rect 3342 2260 3402 2267
rect 4343 1147 4393 1153
rect 4343 1120 4354 1147
rect 4381 1120 4393 1147
rect 4343 1113 4393 1120
rect 3540 954 3580 960
rect 3540 927 3546 954
rect 3573 927 3580 954
rect 3540 920 3580 927
rect 3340 885 3400 892
rect 3340 849 3346 885
rect 3394 849 3400 885
rect 3340 842 3400 849
rect 3341 801 3401 808
rect 3341 765 3347 801
rect 3395 765 3401 801
rect 3341 758 3401 765
rect 3446 736 3489 748
rect 3546 736 3573 920
rect 4354 776 4381 1113
rect 4463 855 4513 860
rect 4783 858 4843 865
rect 4783 855 4788 858
rect 4463 854 4788 855
rect 4463 827 4474 854
rect 4501 827 4788 854
rect 4463 825 4788 827
rect 4463 820 4513 825
rect 4783 822 4788 825
rect 4836 822 4843 858
rect 3446 709 3453 736
rect 3480 709 3573 736
rect 3941 749 4381 776
rect 3446 700 3489 709
rect 3941 493 3968 749
rect 4474 720 4501 820
rect 4783 815 4843 822
rect 3407 466 3968 493
rect 3996 693 4501 720
rect 3407 430 3434 466
rect 3996 430 4023 693
rect 3396 424 3446 430
rect 3396 397 3407 424
rect 3434 397 3446 424
rect 3396 390 3446 397
rect 3985 424 4035 430
rect 3985 397 3996 424
rect 4023 397 4035 424
rect 3985 390 4035 397
rect 3396 268 4759 286
rect 3396 189 3537 268
rect 3659 189 3837 268
rect 3959 189 4137 268
rect 4259 189 4437 268
rect 4559 189 4759 268
rect 3396 177 4759 189
<< via1 >>
rect 3537 2379 3659 2458
rect 3837 2379 3959 2458
rect 4137 2379 4259 2458
rect 4437 2379 4559 2458
rect 3348 2267 3396 2303
rect 3346 849 3394 885
rect 3347 765 3395 801
rect 4788 822 4836 858
rect 3537 189 3659 268
rect 3837 189 3959 268
rect 4137 189 4259 268
rect 4437 189 4559 268
<< metal2 >>
rect 3399 2458 4760 2477
rect 3399 2379 3537 2458
rect 3659 2379 3837 2458
rect 3959 2379 4137 2458
rect 4259 2379 4437 2458
rect 4559 2379 4760 2458
rect 3399 2366 4760 2379
rect 3342 2303 3402 2310
rect 3342 2267 3348 2303
rect 3396 2267 3402 2303
rect 3342 2260 3402 2267
rect 3340 885 3400 892
rect 3340 849 3346 885
rect 3394 849 3400 885
rect 3340 842 3400 849
rect 4783 858 4843 865
rect 4783 822 4788 858
rect 4836 822 4843 858
rect 4783 815 4843 822
rect 3341 801 3401 808
rect 3341 765 3347 801
rect 3395 765 3401 801
rect 3341 758 3401 765
rect 3395 268 4760 286
rect 3395 189 3537 268
rect 3659 189 3837 268
rect 3959 189 4137 268
rect 4259 189 4437 268
rect 4559 189 4760 268
rect 3395 176 4760 189
<< via2 >>
rect 3537 2379 3659 2458
rect 3837 2379 3959 2458
rect 4137 2379 4259 2458
rect 4437 2379 4559 2458
rect 3348 2267 3396 2303
rect 3346 849 3394 885
rect 4788 822 4836 858
rect 3347 765 3395 801
rect 3537 189 3659 268
rect 3837 189 3959 268
rect 4137 189 4259 268
rect 4437 189 4559 268
<< metal3 >>
rect 3399 2458 4760 2477
rect 3399 2379 3537 2458
rect 3659 2379 3837 2458
rect 3959 2379 4137 2458
rect 4259 2379 4437 2458
rect 4559 2379 4760 2458
rect 3399 2366 4760 2379
rect 3342 2303 3402 2310
rect 3342 2267 3348 2303
rect 3396 2267 3402 2303
rect 3342 2260 3402 2267
rect 3340 885 3400 892
rect 3340 849 3346 885
rect 3394 849 3400 885
rect 3340 842 3400 849
rect 4783 858 4843 865
rect 4783 822 4788 858
rect 4836 822 4843 858
rect 4783 815 4843 822
rect 3341 801 3401 808
rect 3341 765 3347 801
rect 3395 765 3401 801
rect 3341 758 3401 765
rect 3395 268 4760 286
rect 3395 189 3537 268
rect 3659 189 3837 268
rect 3959 189 4137 268
rect 4259 189 4437 268
rect 4559 189 4760 268
rect 3395 176 4760 189
<< via3 >>
rect 3348 2267 3396 2303
rect 3346 849 3394 885
rect 4788 822 4836 858
rect 3347 765 3395 801
<< metal4 >>
rect 3342 2303 3402 2310
rect 3342 2267 3348 2303
rect 3396 2267 3402 2303
rect 3342 2260 3402 2267
rect 3340 885 3400 892
rect 3340 849 3346 885
rect 3394 849 3400 885
rect 3340 842 3400 849
rect 4783 858 4843 865
rect 4783 822 4788 858
rect 4836 822 4843 858
rect 4783 815 4843 822
rect 3341 801 3401 808
rect 3341 765 3347 801
rect 3395 765 3401 801
rect 3341 758 3401 765
<< labels >>
flabel metal3 3967 179 4121 278 0 FreeSans 240 0 0 0 VSS
port 5 nsew
flabel metal3 3984 2368 4128 2470 0 FreeSans 240 0 0 0 VDD
port 4 nsew
flabel metal4 3346 764 3396 801 0 FreeSans 240 0 0 0 Inn
port 2 nsew
flabel metal4 3346 849 3394 885 0 FreeSans 240 0 0 0 Inp
port 1 nsew
flabel metal4 3347 2263 3398 2305 0 FreeSans 240 0 0 0 Ib
port 6 nsew
flabel metal4 4787 822 4835 858 0 FreeSans 160 0 0 0 vout
port 3 nsew
<< end >>
