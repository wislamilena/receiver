magic
tech sky130A
magscale 1 2
timestamp 1647797958
<< pwell >>
rect -45690 -11880 -45550 -7380
<< nmos >>
rect -45860 -11880 -45830 -7380
<< ndiff >>
rect -46000 -7459 -45860 -7380
rect -46000 -7493 -45943 -7459
rect -45909 -7493 -45860 -7459
rect -46000 -7527 -45860 -7493
rect -46000 -7561 -45943 -7527
rect -45909 -7561 -45860 -7527
rect -46000 -8298 -45860 -7561
rect -46000 -8332 -45941 -8298
rect -45907 -8332 -45860 -8298
rect -46000 -8366 -45860 -8332
rect -46000 -8400 -45941 -8366
rect -45907 -8400 -45860 -8366
rect -46000 -8999 -45860 -8400
rect -46000 -9033 -45941 -8999
rect -45907 -9033 -45860 -8999
rect -46000 -9067 -45860 -9033
rect -46000 -9101 -45941 -9067
rect -45907 -9101 -45860 -9067
rect -46000 -10299 -45860 -9101
rect -46000 -10333 -45941 -10299
rect -45907 -10333 -45860 -10299
rect -46000 -10367 -45860 -10333
rect -46000 -10401 -45941 -10367
rect -45907 -10401 -45860 -10367
rect -46000 -11599 -45860 -10401
rect -46000 -11633 -45941 -11599
rect -45907 -11633 -45860 -11599
rect -46000 -11667 -45860 -11633
rect -46000 -11701 -45941 -11667
rect -45907 -11701 -45860 -11667
rect -46000 -11880 -45860 -11701
rect -45830 -7453 -45690 -7380
rect -45830 -7487 -45751 -7453
rect -45717 -7487 -45690 -7453
rect -45830 -7521 -45690 -7487
rect -45830 -7555 -45751 -7521
rect -45717 -7555 -45690 -7521
rect -45830 -7899 -45690 -7555
rect -45830 -7933 -45753 -7899
rect -45719 -7933 -45690 -7899
rect -45830 -7967 -45690 -7933
rect -45830 -8001 -45753 -7967
rect -45719 -8001 -45690 -7967
rect -45830 -8405 -45690 -8001
rect -45830 -8439 -45749 -8405
rect -45715 -8439 -45690 -8405
rect -45830 -8473 -45690 -8439
rect -45830 -8507 -45749 -8473
rect -45715 -8507 -45690 -8473
rect -45830 -9193 -45690 -8507
rect -45830 -9227 -45761 -9193
rect -45727 -9227 -45690 -9193
rect -45830 -9261 -45690 -9227
rect -45830 -9295 -45761 -9261
rect -45727 -9295 -45690 -9261
rect -45830 -9799 -45690 -9295
rect -45830 -9833 -45755 -9799
rect -45721 -9833 -45690 -9799
rect -45830 -9867 -45690 -9833
rect -45830 -9901 -45755 -9867
rect -45721 -9901 -45690 -9867
rect -45830 -10405 -45690 -9901
rect -45830 -10439 -45749 -10405
rect -45715 -10439 -45690 -10405
rect -45830 -10473 -45690 -10439
rect -45830 -10507 -45749 -10473
rect -45715 -10507 -45690 -10473
rect -45830 -11603 -45690 -10507
rect -45830 -11637 -45751 -11603
rect -45717 -11637 -45690 -11603
rect -45830 -11671 -45690 -11637
rect -45830 -11705 -45751 -11671
rect -45717 -11705 -45690 -11671
rect -45830 -11880 -45690 -11705
<< ndiffc >>
rect -45943 -7493 -45909 -7459
rect -45943 -7561 -45909 -7527
rect -45941 -8332 -45907 -8298
rect -45941 -8400 -45907 -8366
rect -45941 -9033 -45907 -8999
rect -45941 -9101 -45907 -9067
rect -45941 -10333 -45907 -10299
rect -45941 -10401 -45907 -10367
rect -45941 -11633 -45907 -11599
rect -45941 -11701 -45907 -11667
rect -45751 -7487 -45717 -7453
rect -45751 -7555 -45717 -7521
rect -45753 -7933 -45719 -7899
rect -45753 -8001 -45719 -7967
rect -45749 -8439 -45715 -8405
rect -45749 -8507 -45715 -8473
rect -45761 -9227 -45727 -9193
rect -45761 -9295 -45727 -9261
rect -45755 -9833 -45721 -9799
rect -45755 -9901 -45721 -9867
rect -45749 -10439 -45715 -10405
rect -45749 -10507 -45715 -10473
rect -45751 -11637 -45717 -11603
rect -45751 -11705 -45717 -11671
<< psubdiff >>
rect -45690 -7459 -45550 -7380
rect -45690 -7493 -45657 -7459
rect -45623 -7493 -45550 -7459
rect -45690 -7527 -45550 -7493
rect -45690 -7561 -45657 -7527
rect -45623 -7561 -45550 -7527
rect -45690 -7899 -45550 -7561
rect -45690 -7933 -45657 -7899
rect -45623 -7933 -45550 -7899
rect -45690 -7967 -45550 -7933
rect -45690 -8001 -45657 -7967
rect -45623 -8001 -45550 -7967
rect -45690 -8409 -45550 -8001
rect -45690 -8443 -45653 -8409
rect -45619 -8443 -45550 -8409
rect -45690 -8477 -45550 -8443
rect -45690 -8511 -45653 -8477
rect -45619 -8511 -45550 -8477
rect -45690 -9199 -45550 -8511
rect -45690 -9233 -45655 -9199
rect -45621 -9233 -45550 -9199
rect -45690 -9267 -45550 -9233
rect -45690 -9301 -45655 -9267
rect -45621 -9301 -45550 -9267
rect -45690 -9799 -45550 -9301
rect -45690 -9833 -45657 -9799
rect -45623 -9833 -45550 -9799
rect -45690 -9867 -45550 -9833
rect -45690 -9901 -45657 -9867
rect -45623 -9901 -45550 -9867
rect -45690 -10409 -45550 -9901
rect -45690 -10443 -45653 -10409
rect -45619 -10443 -45550 -10409
rect -45690 -10477 -45550 -10443
rect -45690 -10511 -45653 -10477
rect -45619 -10511 -45550 -10477
rect -45690 -11599 -45550 -10511
rect -45690 -11633 -45657 -11599
rect -45623 -11633 -45550 -11599
rect -45690 -11667 -45550 -11633
rect -45690 -11701 -45657 -11667
rect -45623 -11701 -45550 -11667
rect -45690 -11880 -45550 -11701
<< psubdiffcont >>
rect -45657 -7493 -45623 -7459
rect -45657 -7561 -45623 -7527
rect -45657 -7933 -45623 -7899
rect -45657 -8001 -45623 -7967
rect -45653 -8443 -45619 -8409
rect -45653 -8511 -45619 -8477
rect -45655 -9233 -45621 -9199
rect -45655 -9301 -45621 -9267
rect -45657 -9833 -45623 -9799
rect -45657 -9901 -45623 -9867
rect -45653 -10443 -45619 -10409
rect -45653 -10511 -45619 -10477
rect -45657 -11633 -45623 -11599
rect -45657 -11701 -45623 -11667
<< poly >>
rect -45860 -7380 -45830 -7280
rect -45860 -11996 -45830 -11880
rect -45934 -12013 -45754 -11996
rect -45934 -12047 -45862 -12013
rect -45828 -12047 -45754 -12013
rect -45934 -12080 -45754 -12047
<< polycont >>
rect -45862 -12047 -45828 -12013
<< locali >>
rect -52120 -3207 -39006 -2992
rect -52120 -3745 -50981 -3207
rect -50011 -3745 -47981 -3207
rect -47011 -3745 -44981 -3207
rect -44011 -3227 -39006 -3207
rect -44011 -3745 -40771 -3227
rect -52120 -3765 -40771 -3745
rect -40233 -3765 -39006 -3227
rect -52120 -4028 -39006 -3765
rect -46010 -5492 -45840 -5458
rect -46010 -5526 -45945 -5492
rect -45911 -5526 -45840 -5492
rect -46010 -5570 -45840 -5526
rect -45970 -7459 -45886 -5570
rect -45730 -7420 -45650 -4028
rect -45970 -7493 -45943 -7459
rect -45909 -7493 -45886 -7459
rect -45970 -7527 -45886 -7493
rect -45970 -7561 -45943 -7527
rect -45909 -7561 -45886 -7527
rect -45970 -7590 -45886 -7561
rect -45780 -7453 -45586 -7420
rect -45780 -7487 -45751 -7453
rect -45717 -7459 -45586 -7453
rect -45717 -7487 -45657 -7459
rect -45780 -7493 -45657 -7487
rect -45623 -7493 -45586 -7459
rect -45780 -7521 -45586 -7493
rect -45780 -7555 -45751 -7521
rect -45717 -7527 -45586 -7521
rect -45717 -7555 -45657 -7527
rect -45780 -7561 -45657 -7555
rect -45623 -7561 -45586 -7527
rect -45780 -7590 -45586 -7561
rect -45784 -7899 -45590 -7858
rect -45784 -7933 -45753 -7899
rect -45719 -7933 -45657 -7899
rect -45623 -7933 -45590 -7899
rect -45784 -7967 -45590 -7933
rect -45784 -8001 -45753 -7967
rect -45719 -8001 -45657 -7967
rect -45623 -8001 -45590 -7967
rect -45784 -8028 -45590 -8001
rect -45970 -8298 -45876 -8270
rect -45970 -8332 -45941 -8298
rect -45907 -8332 -45876 -8298
rect -45970 -8366 -45876 -8332
rect -45970 -8400 -45941 -8366
rect -45907 -8400 -45876 -8366
rect -45970 -8430 -45876 -8400
rect -45780 -8405 -45588 -8370
rect -45780 -8439 -45749 -8405
rect -45715 -8409 -45588 -8405
rect -45715 -8439 -45653 -8409
rect -45780 -8443 -45653 -8439
rect -45619 -8443 -45588 -8409
rect -45780 -8473 -45588 -8443
rect -45780 -8507 -45749 -8473
rect -45715 -8477 -45588 -8473
rect -45715 -8507 -45653 -8477
rect -45780 -8511 -45653 -8507
rect -45619 -8511 -45588 -8477
rect -45780 -8540 -45588 -8511
rect -45970 -8999 -45876 -8970
rect -45970 -9033 -45941 -8999
rect -45907 -9033 -45876 -8999
rect -45970 -9067 -45876 -9033
rect -45970 -9101 -45941 -9067
rect -45907 -9101 -45876 -9067
rect -45970 -9130 -45876 -9101
rect -45790 -9193 -45590 -9160
rect -45790 -9227 -45761 -9193
rect -45727 -9199 -45590 -9193
rect -45727 -9227 -45655 -9199
rect -45790 -9233 -45655 -9227
rect -45621 -9233 -45590 -9199
rect -45790 -9261 -45590 -9233
rect -45790 -9295 -45761 -9261
rect -45727 -9267 -45590 -9261
rect -45727 -9295 -45655 -9267
rect -45790 -9301 -45655 -9295
rect -45621 -9301 -45590 -9267
rect -45790 -9330 -45590 -9301
rect -45784 -9799 -45590 -9758
rect -45784 -9833 -45755 -9799
rect -45721 -9833 -45657 -9799
rect -45623 -9833 -45590 -9799
rect -45784 -9867 -45590 -9833
rect -45784 -9901 -45755 -9867
rect -45721 -9901 -45657 -9867
rect -45623 -9901 -45590 -9867
rect -45784 -9928 -45590 -9901
rect -45970 -10299 -45876 -10270
rect -45970 -10333 -45941 -10299
rect -45907 -10333 -45876 -10299
rect -45970 -10367 -45876 -10333
rect -45970 -10401 -45941 -10367
rect -45907 -10401 -45876 -10367
rect -45970 -10430 -45876 -10401
rect -45780 -10405 -45588 -10370
rect -45780 -10439 -45749 -10405
rect -45715 -10409 -45588 -10405
rect -45715 -10439 -45653 -10409
rect -45780 -10443 -45653 -10439
rect -45619 -10443 -45588 -10409
rect -45780 -10473 -45588 -10443
rect -45780 -10507 -45749 -10473
rect -45715 -10477 -45588 -10473
rect -45715 -10507 -45653 -10477
rect -45780 -10511 -45653 -10507
rect -45619 -10511 -45588 -10477
rect -45780 -10540 -45588 -10511
rect -45970 -11599 -45876 -11570
rect -45970 -11633 -45941 -11599
rect -45907 -11633 -45876 -11599
rect -45970 -11667 -45876 -11633
rect -45970 -11701 -45941 -11667
rect -45907 -11701 -45876 -11667
rect -45970 -11730 -45876 -11701
rect -45780 -11599 -45588 -11570
rect -45780 -11603 -45657 -11599
rect -45780 -11637 -45751 -11603
rect -45717 -11633 -45657 -11603
rect -45623 -11633 -45588 -11599
rect -45717 -11637 -45588 -11633
rect -45780 -11667 -45588 -11637
rect -45780 -11671 -45657 -11667
rect -45780 -11705 -45751 -11671
rect -45717 -11701 -45657 -11671
rect -45623 -11701 -45588 -11667
rect -45717 -11705 -45588 -11701
rect -45780 -11740 -45588 -11705
rect -46122 -12013 -45526 -11996
rect -46122 -12047 -45862 -12013
rect -45828 -12047 -45526 -12013
rect -46122 -26620 -45526 -12047
<< viali >>
rect -50981 -3745 -50011 -3207
rect -47981 -3745 -47011 -3207
rect -44981 -3745 -44011 -3207
rect -40771 -3765 -40233 -3227
rect -45945 -5526 -45911 -5492
<< metal1 >>
rect -52120 -3207 -39006 -2992
rect -52120 -3745 -50981 -3207
rect -50011 -3745 -47981 -3207
rect -47011 -3745 -44981 -3207
rect -44011 -3214 -39006 -3207
rect -44011 -3745 -40784 -3214
rect -52120 -3778 -40784 -3745
rect -40220 -3778 -39006 -3214
rect -52120 -4028 -39006 -3778
rect -46010 -5483 -45840 -5458
rect -46010 -5535 -45954 -5483
rect -45902 -5535 -45840 -5483
rect -44800 -5464 -44680 -5450
rect -44800 -5516 -44768 -5464
rect -44716 -5516 -44680 -5464
rect -44800 -5530 -44680 -5516
rect -46010 -5570 -45840 -5535
rect -44770 -7044 -44700 -5530
rect -44760 -11620 -44710 -11612
rect -44770 -12551 -44700 -11620
rect -44936 -25000 -44534 -12551
rect -42992 -24904 -41392 -24390
rect -42992 -25000 -42484 -24904
rect -44936 -25342 -42484 -25000
rect -44936 -25356 -44534 -25342
rect -42992 -25468 -42484 -25342
rect -41920 -25468 -41392 -24904
rect -42992 -25990 -41392 -25468
<< via1 >>
rect -40784 -3227 -40220 -3214
rect -40784 -3765 -40771 -3227
rect -40771 -3765 -40233 -3227
rect -40233 -3765 -40220 -3227
rect -40784 -3778 -40220 -3765
rect -45954 -5492 -45902 -5483
rect -45954 -5526 -45945 -5492
rect -45945 -5526 -45911 -5492
rect -45911 -5526 -45902 -5492
rect -45954 -5535 -45902 -5526
rect -44768 -5516 -44716 -5464
rect -42484 -25468 -41920 -24904
<< metal2 >>
rect -40996 -3214 -39992 -3004
rect -40996 -3778 -40784 -3214
rect -40220 -3778 -39992 -3214
rect -40996 -4008 -39992 -3778
rect -46010 -5481 -45840 -5458
rect -46010 -5537 -45956 -5481
rect -45900 -5537 -45840 -5481
rect -44800 -5462 -44680 -5450
rect -44800 -5518 -44770 -5462
rect -44714 -5518 -44680 -5462
rect -44800 -5530 -44680 -5518
rect -46010 -5570 -45840 -5537
rect -42992 -24904 -41392 -24390
rect -42992 -25468 -42484 -24904
rect -41920 -25468 -41392 -24904
rect -42992 -25990 -41392 -25468
<< via2 >>
rect -40770 -3764 -40234 -3228
rect -45956 -5483 -45900 -5481
rect -45956 -5535 -45954 -5483
rect -45954 -5535 -45902 -5483
rect -45902 -5535 -45900 -5483
rect -45956 -5537 -45900 -5535
rect -44770 -5464 -44714 -5462
rect -44770 -5516 -44768 -5464
rect -44768 -5516 -44716 -5464
rect -44716 -5516 -44714 -5464
rect -44770 -5518 -44714 -5516
rect -42470 -25454 -41934 -24918
<< metal3 >>
rect -41006 -3228 -40002 -3000
rect -41006 -3764 -40770 -3228
rect -40234 -3764 -40002 -3228
rect -41006 -4800 -40002 -3764
rect -47686 -5000 -44398 -4998
rect -49400 -5002 -44398 -5000
rect -49400 -5462 -44392 -5002
rect -41004 -5400 -39998 -4800
rect -49400 -5481 -44770 -5462
rect -49400 -5537 -45956 -5481
rect -45900 -5518 -44770 -5481
rect -44714 -5518 -44392 -5462
rect -45900 -5537 -44392 -5518
rect -49400 -5600 -44392 -5537
rect -49400 -5602 -44398 -5600
rect -49400 -6208 -48400 -5602
rect -41002 -6188 -40002 -5400
rect -64974 -23788 -47386 -6208
rect -43100 -23782 -25500 -6188
rect -42992 -24914 -41392 -24390
rect -42992 -25458 -42474 -24914
rect -41930 -25458 -41392 -24914
rect -42992 -25990 -41392 -25458
<< via3 >>
rect -42474 -24918 -41930 -24914
rect -42474 -25454 -42470 -24918
rect -42470 -25454 -41934 -24918
rect -41934 -25454 -41930 -24918
rect -42474 -25458 -41930 -25454
<< mimcap >>
rect -64884 -16971 -47484 -6308
rect -64884 -19995 -62437 -16971
rect -58133 -19995 -47484 -16971
rect -64884 -23708 -47484 -19995
rect -43000 -16629 -25600 -6276
rect -43000 -19653 -40023 -16629
rect -35719 -19653 -25600 -16629
rect -43000 -23676 -25600 -19653
<< mimcapcontact >>
rect -62437 -19995 -58133 -16971
rect -40023 -19653 -35719 -16629
<< metal4 >>
rect -63034 -16971 -57576 -16188
rect -63034 -19995 -62437 -16971
rect -58133 -19995 -57576 -16971
rect -63034 -26814 -57576 -19995
rect -40492 -16629 -35034 -15568
rect -40492 -19653 -40023 -16629
rect -35719 -19653 -35034 -16629
rect -42992 -24914 -41392 -24390
rect -42992 -25458 -42474 -24914
rect -41930 -25008 -41392 -24914
rect -40492 -25008 -35034 -19653
rect -41930 -25350 -35034 -25008
rect -41930 -25458 -41392 -25350
rect -42992 -25990 -41392 -25458
rect -40492 -26942 -35034 -25350
use sky130_fd_pr__res_xhigh_po_0p35_HDW2JU  R
timestamp 1647797958
transform 1 0 -44735 0 1 -9330
box -35 -2292 35 2292
<< labels >>
flabel metal3 s -49252 -5534 -48136 -5026 0 FreeSans 1250 0 0 0 bot_cin
rlabel metal4 s -63034 -25264 -63034 -25264 4 din
port 1 nsew
rlabel locali s -45852 -26620 -45852 -26620 4 db
port 2 nsew
rlabel metal4 s -35040 -25176 -35040 -25176 4 do
port 3 nsew
rlabel metal1 s -52114 -3556 -52114 -3556 4 GND
port 4 nsew
<< end >>
