magic
tech sky130A
magscale 1 2
timestamp 1647797958
<< xpolycontact >>
rect -35 1860 35 2292
rect -35 -2292 35 -1860
<< xpolyres >>
rect -35 -1860 35 1860
<< viali >>
rect -17 2238 17 2272
rect -17 2166 17 2200
rect -17 2094 17 2128
rect -17 2022 17 2056
rect -17 1950 17 1984
rect -17 1878 17 1912
rect -17 -1913 17 -1879
rect -17 -1985 17 -1951
rect -17 -2057 17 -2023
rect -17 -2129 17 -2095
rect -17 -2201 17 -2167
rect -17 -2273 17 -2239
<< metal1 >>
rect -25 2272 25 2286
rect -25 2238 -17 2272
rect 17 2238 25 2272
rect -25 2200 25 2238
rect -25 2166 -17 2200
rect 17 2166 25 2200
rect -25 2128 25 2166
rect -25 2094 -17 2128
rect 17 2094 25 2128
rect -25 2056 25 2094
rect -25 2022 -17 2056
rect 17 2022 25 2056
rect -25 1984 25 2022
rect -25 1950 -17 1984
rect 17 1950 25 1984
rect -25 1912 25 1950
rect -25 1878 -17 1912
rect 17 1878 25 1912
rect -25 1865 25 1878
rect -25 -1879 25 -1865
rect -25 -1913 -17 -1879
rect 17 -1913 25 -1879
rect -25 -1951 25 -1913
rect -25 -1985 -17 -1951
rect 17 -1985 25 -1951
rect -25 -2023 25 -1985
rect -25 -2057 -17 -2023
rect 17 -2057 25 -2023
rect -25 -2095 25 -2057
rect -25 -2129 -17 -2095
rect 17 -2129 25 -2095
rect -25 -2167 25 -2129
rect -25 -2201 -17 -2167
rect 17 -2201 25 -2167
rect -25 -2239 25 -2201
rect -25 -2273 -17 -2239
rect 17 -2273 25 -2239
rect -25 -2286 25 -2273
<< end >>
