* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p35_HDW2JU a_n35_1860# a_n35_n2292# VSUBS
X0 a_n35_n2292# a_n35_1860# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=1.86e+07u
C0 a_n35_n2292# VSUBS 0.55fF
C1 a_n35_1860# VSUBS 0.55fF
.ends

.subckt detV2 din db do GND
XR a_n46000_n11880# do GND sky130_fd_pr__res_xhigh_po_0p35_HDW2JU
X0 din a_n46000_n11880# sky130_fd_pr__cap_mim_m3_1 l=8.7e+07u w=8.7e+07u
X1 do GND sky130_fd_pr__cap_mim_m3_1 l=8.7e+07u w=8.7e+07u
X2 GND db a_n46000_n11880# GND sky130_fd_pr__nfet_01v8 w=2.25e+07u l=150000u
C0 db a_n46000_n11880# 0.01fF
C1 din a_n46000_n11880# 95.06fF
C2 din GND 5.50fF
C3 db GND 16.77fF
C4 do GND 125.35fF
C5 a_n46000_n11880# GND 112.58fF
.ends

.subckt user_analog_project_wrapper
XdetV2_0 io_analog[2] detV2_0/db io_analog[3] vssa1 detV2
C0 user_analog_project_wrapper_empty_0/io_clamp_high[1] user_analog_project_wrapper_empty_0/io_analog[5] 0.53fF
C1 user_analog_project_wrapper_empty_0/io_clamp_high[0] user_analog_project_wrapper_empty_0/io_clamp_low[0] 0.53fF
C2 user_analog_project_wrapper_empty_0/io_clamp_high[1] user_analog_project_wrapper_empty_0/io_clamp_low[1] 0.53fF
C3 io_analog[2] detV2_0/db 10.68fF
C4 user_analog_project_wrapper_empty_0/io_analog[5] user_analog_project_wrapper_empty_0/io_clamp_low[1] 0.53fF
C5 user_analog_project_wrapper_empty_0/io_clamp_high[2] user_analog_project_wrapper_empty_0/io_analog[6] 0.53fF
C6 user_analog_project_wrapper_empty_0/io_clamp_high[0] user_analog_project_wrapper_empty_0/io_analog[4] 0.53fF
C7 user_analog_project_wrapper_empty_0/io_clamp_low[2] user_analog_project_wrapper_empty_0/io_analog[6] 0.53fF
C8 user_analog_project_wrapper_empty_0/io_clamp_low[2] user_analog_project_wrapper_empty_0/io_clamp_high[2] 0.53fF
C9 user_analog_project_wrapper_empty_0/io_analog[4] user_analog_project_wrapper_empty_0/io_clamp_low[0] 0.53fF
C10 io_analog[2] vssa1 154.95fF
C11 detV2_0/db vssa1 230.22fF
C12 io_analog[3] vssa1 199.92fF
C13 detV2_0/a_n46000_n11880# vssa1 112.58fF
C14 user_analog_project_wrapper_empty_0/io_analog[4] vssa1 25.05fF
C15 user_analog_project_wrapper_empty_0/io_analog[5] vssa1 25.05fF
C16 user_analog_project_wrapper_empty_0/io_analog[6] vssa1 25.05fF
C17 user_analog_project_wrapper_empty_0/io_in_3v3[0] vssa1 0.61fF
C18 user_analog_project_wrapper_empty_0/io_oeb[26] vssa1 0.61fF
C19 user_analog_project_wrapper_empty_0/io_in[0] vssa1 0.61fF
C20 user_analog_project_wrapper_empty_0/io_out[26] vssa1 0.61fF
C21 user_analog_project_wrapper_empty_0/io_out[0] vssa1 0.61fF
C22 user_analog_project_wrapper_empty_0/io_in[26] vssa1 0.61fF
C23 user_analog_project_wrapper_empty_0/io_oeb[0] vssa1 0.61fF
C24 user_analog_project_wrapper_empty_0/io_in_3v3[26] vssa1 0.61fF
C25 user_analog_project_wrapper_empty_0/io_in_3v3[1] vssa1 0.61fF
C26 user_analog_project_wrapper_empty_0/io_oeb[25] vssa1 0.61fF
C27 user_analog_project_wrapper_empty_0/io_in[1] vssa1 0.61fF
C28 user_analog_project_wrapper_empty_0/io_out[25] vssa1 0.61fF
C29 user_analog_project_wrapper_empty_0/io_out[1] vssa1 0.61fF
C30 user_analog_project_wrapper_empty_0/io_in[25] vssa1 0.61fF
C31 user_analog_project_wrapper_empty_0/io_oeb[1] vssa1 0.61fF
C32 user_analog_project_wrapper_empty_0/io_in_3v3[25] vssa1 0.61fF
C33 user_analog_project_wrapper_empty_0/io_in_3v3[2] vssa1 0.61fF
C34 user_analog_project_wrapper_empty_0/io_oeb[24] vssa1 0.61fF
C35 user_analog_project_wrapper_empty_0/io_in[2] vssa1 0.61fF
C36 user_analog_project_wrapper_empty_0/io_out[24] vssa1 0.61fF
C37 user_analog_project_wrapper_empty_0/io_out[2] vssa1 0.61fF
C38 user_analog_project_wrapper_empty_0/io_in[24] vssa1 0.61fF
C39 user_analog_project_wrapper_empty_0/io_oeb[2] vssa1 0.61fF
C40 user_analog_project_wrapper_empty_0/io_in_3v3[24] vssa1 0.61fF
C41 user_analog_project_wrapper_empty_0/io_in_3v3[3] vssa1 0.61fF
C42 user_analog_project_wrapper_empty_0/gpio_noesd[17] vssa1 0.61fF
C43 user_analog_project_wrapper_empty_0/io_in[3] vssa1 0.61fF
C44 user_analog_project_wrapper_empty_0/gpio_analog[17] vssa1 0.61fF
C45 user_analog_project_wrapper_empty_0/io_out[3] vssa1 0.61fF
C46 user_analog_project_wrapper_empty_0/io_oeb[3] vssa1 0.61fF
C47 user_analog_project_wrapper_empty_0/io_in_3v3[4] vssa1 0.61fF
C48 user_analog_project_wrapper_empty_0/io_in[4] vssa1 0.61fF
C49 user_analog_project_wrapper_empty_0/io_out[4] vssa1 0.61fF
C50 user_analog_project_wrapper_empty_0/io_oeb[4] vssa1 0.61fF
C51 user_analog_project_wrapper_empty_0/io_oeb[23] vssa1 0.61fF
C52 user_analog_project_wrapper_empty_0/io_out[23] vssa1 0.61fF
C53 user_analog_project_wrapper_empty_0/io_in[23] vssa1 0.61fF
C54 user_analog_project_wrapper_empty_0/io_in_3v3[23] vssa1 0.61fF
C55 user_analog_project_wrapper_empty_0/gpio_noesd[16] vssa1 0.61fF
C56 user_analog_project_wrapper_empty_0/gpio_analog[16] vssa1 0.61fF
C57 user_analog_project_wrapper_empty_0/io_in_3v3[5] vssa1 0.61fF
C58 user_analog_project_wrapper_empty_0/io_in[5] vssa1 0.61fF
C59 user_analog_project_wrapper_empty_0/io_out[5] vssa1 0.61fF
C60 user_analog_project_wrapper_empty_0/io_oeb[5] vssa1 0.61fF
C61 user_analog_project_wrapper_empty_0/io_oeb[22] vssa1 0.61fF
C62 user_analog_project_wrapper_empty_0/io_out[22] vssa1 0.61fF
C63 user_analog_project_wrapper_empty_0/io_in[22] vssa1 0.61fF
C64 user_analog_project_wrapper_empty_0/io_in_3v3[22] vssa1 0.61fF
C65 user_analog_project_wrapper_empty_0/gpio_noesd[15] vssa1 0.61fF
C66 user_analog_project_wrapper_empty_0/gpio_analog[15] vssa1 0.61fF
C67 user_analog_project_wrapper_empty_0/io_in_3v3[6] vssa1 0.61fF
C68 user_analog_project_wrapper_empty_0/io_in[6] vssa1 0.61fF
C69 user_analog_project_wrapper_empty_0/io_out[6] vssa1 0.61fF
C70 user_analog_project_wrapper_empty_0/io_oeb[6] vssa1 0.61fF
C71 user_analog_project_wrapper_empty_0/io_oeb[21] vssa1 0.61fF
C72 user_analog_project_wrapper_empty_0/io_out[21] vssa1 0.61fF
C73 user_analog_project_wrapper_empty_0/io_in[21] vssa1 0.61fF
C74 user_analog_project_wrapper_empty_0/io_in_3v3[21] vssa1 0.61fF
C75 user_analog_project_wrapper_empty_0/gpio_noesd[14] vssa1 0.61fF
C76 user_analog_project_wrapper_empty_0/gpio_analog[14] vssa1 0.61fF
C77 user_analog_project_wrapper_empty_0/vssd2 vssa1 13.04fF
C78 user_analog_project_wrapper_empty_0/vssd1 vssa1 13.04fF
C79 user_analog_project_wrapper_empty_0/vdda2 vssa1 13.04fF
C80 user_analog_project_wrapper_empty_0/vdda1 vssa1 26.08fF
C81 user_analog_project_wrapper_empty_0/io_oeb[20] vssa1 0.61fF
C82 user_analog_project_wrapper_empty_0/io_out[20] vssa1 0.61fF
C83 user_analog_project_wrapper_empty_0/io_in[20] vssa1 0.61fF
C84 user_analog_project_wrapper_empty_0/io_in_3v3[20] vssa1 0.61fF
C85 user_analog_project_wrapper_empty_0/gpio_noesd[13] vssa1 0.61fF
C86 user_analog_project_wrapper_empty_0/gpio_analog[13] vssa1 0.61fF
C87 user_analog_project_wrapper_empty_0/gpio_analog[0] vssa1 0.61fF
C88 user_analog_project_wrapper_empty_0/gpio_noesd[0] vssa1 0.61fF
C89 user_analog_project_wrapper_empty_0/io_in_3v3[7] vssa1 0.61fF
C90 user_analog_project_wrapper_empty_0/io_in[7] vssa1 0.61fF
C91 user_analog_project_wrapper_empty_0/io_out[7] vssa1 0.61fF
C92 user_analog_project_wrapper_empty_0/io_oeb[7] vssa1 0.61fF
C93 user_analog_project_wrapper_empty_0/io_oeb[19] vssa1 0.61fF
C94 user_analog_project_wrapper_empty_0/io_out[19] vssa1 0.61fF
C95 user_analog_project_wrapper_empty_0/io_in[19] vssa1 0.61fF
C96 user_analog_project_wrapper_empty_0/io_in_3v3[19] vssa1 0.61fF
C97 user_analog_project_wrapper_empty_0/gpio_noesd[12] vssa1 0.61fF
C98 user_analog_project_wrapper_empty_0/gpio_analog[12] vssa1 0.61fF
C99 user_analog_project_wrapper_empty_0/gpio_analog[1] vssa1 0.61fF
C100 user_analog_project_wrapper_empty_0/gpio_noesd[1] vssa1 0.61fF
C101 user_analog_project_wrapper_empty_0/io_in_3v3[8] vssa1 0.61fF
C102 user_analog_project_wrapper_empty_0/io_in[8] vssa1 0.61fF
C103 user_analog_project_wrapper_empty_0/io_out[8] vssa1 0.61fF
C104 user_analog_project_wrapper_empty_0/io_oeb[8] vssa1 0.61fF
C105 user_analog_project_wrapper_empty_0/io_oeb[18] vssa1 0.61fF
C106 user_analog_project_wrapper_empty_0/io_out[18] vssa1 0.61fF
C107 user_analog_project_wrapper_empty_0/io_in[18] vssa1 0.61fF
C108 user_analog_project_wrapper_empty_0/io_in_3v3[18] vssa1 0.61fF
C109 user_analog_project_wrapper_empty_0/gpio_noesd[11] vssa1 0.61fF
C110 user_analog_project_wrapper_empty_0/gpio_analog[11] vssa1 0.61fF
C111 user_analog_project_wrapper_empty_0/gpio_analog[2] vssa1 0.61fF
C112 user_analog_project_wrapper_empty_0/gpio_noesd[2] vssa1 0.61fF
C113 user_analog_project_wrapper_empty_0/io_in_3v3[9] vssa1 0.61fF
C114 user_analog_project_wrapper_empty_0/io_in[9] vssa1 0.61fF
C115 user_analog_project_wrapper_empty_0/io_out[9] vssa1 0.61fF
C116 user_analog_project_wrapper_empty_0/io_oeb[9] vssa1 0.61fF
C117 user_analog_project_wrapper_empty_0/io_oeb[17] vssa1 0.61fF
C118 user_analog_project_wrapper_empty_0/io_out[17] vssa1 0.61fF
C119 user_analog_project_wrapper_empty_0/io_in[17] vssa1 0.61fF
C120 user_analog_project_wrapper_empty_0/io_in_3v3[17] vssa1 0.61fF
C121 user_analog_project_wrapper_empty_0/gpio_noesd[10] vssa1 0.61fF
C122 user_analog_project_wrapper_empty_0/gpio_analog[10] vssa1 0.61fF
C123 user_analog_project_wrapper_empty_0/gpio_analog[3] vssa1 0.61fF
C124 user_analog_project_wrapper_empty_0/gpio_noesd[3] vssa1 0.61fF
C125 user_analog_project_wrapper_empty_0/io_in_3v3[10] vssa1 0.61fF
C126 user_analog_project_wrapper_empty_0/io_in[10] vssa1 0.61fF
C127 user_analog_project_wrapper_empty_0/io_out[10] vssa1 0.61fF
C128 user_analog_project_wrapper_empty_0/io_oeb[10] vssa1 0.61fF
C129 user_analog_project_wrapper_empty_0/io_oeb[16] vssa1 0.61fF
C130 user_analog_project_wrapper_empty_0/io_out[16] vssa1 0.61fF
C131 user_analog_project_wrapper_empty_0/io_in[16] vssa1 0.61fF
C132 user_analog_project_wrapper_empty_0/io_in_3v3[16] vssa1 0.61fF
C133 user_analog_project_wrapper_empty_0/gpio_noesd[9] vssa1 0.61fF
C134 user_analog_project_wrapper_empty_0/gpio_analog[9] vssa1 0.61fF
C135 user_analog_project_wrapper_empty_0/gpio_analog[4] vssa1 0.61fF
C136 user_analog_project_wrapper_empty_0/gpio_noesd[4] vssa1 0.61fF
C137 user_analog_project_wrapper_empty_0/io_in_3v3[11] vssa1 0.61fF
C138 user_analog_project_wrapper_empty_0/io_in[11] vssa1 0.61fF
C139 user_analog_project_wrapper_empty_0/io_out[11] vssa1 0.61fF
C140 user_analog_project_wrapper_empty_0/io_oeb[11] vssa1 0.61fF
C141 user_analog_project_wrapper_empty_0/io_oeb[15] vssa1 0.61fF
C142 user_analog_project_wrapper_empty_0/io_out[15] vssa1 0.61fF
C143 user_analog_project_wrapper_empty_0/io_in[15] vssa1 0.61fF
C144 user_analog_project_wrapper_empty_0/io_in_3v3[15] vssa1 0.61fF
C145 user_analog_project_wrapper_empty_0/gpio_noesd[8] vssa1 0.61fF
C146 user_analog_project_wrapper_empty_0/gpio_analog[8] vssa1 0.61fF
C147 user_analog_project_wrapper_empty_0/gpio_analog[5] vssa1 0.61fF
C148 user_analog_project_wrapper_empty_0/gpio_noesd[5] vssa1 0.61fF
C149 user_analog_project_wrapper_empty_0/io_in_3v3[12] vssa1 0.61fF
C150 user_analog_project_wrapper_empty_0/io_in[12] vssa1 0.61fF
C151 user_analog_project_wrapper_empty_0/io_out[12] vssa1 0.61fF
C152 user_analog_project_wrapper_empty_0/io_oeb[12] vssa1 0.61fF
C153 user_analog_project_wrapper_empty_0/io_oeb[14] vssa1 0.61fF
C154 user_analog_project_wrapper_empty_0/io_out[14] vssa1 0.61fF
C155 user_analog_project_wrapper_empty_0/io_in[14] vssa1 0.61fF
C156 user_analog_project_wrapper_empty_0/io_in_3v3[14] vssa1 0.61fF
C157 user_analog_project_wrapper_empty_0/gpio_noesd[7] vssa1 0.61fF
C158 user_analog_project_wrapper_empty_0/gpio_analog[7] vssa1 0.61fF
C159 user_analog_project_wrapper_empty_0/vssa2 vssa1 13.04fF
C160 user_analog_project_wrapper_empty_0/gpio_analog[6] vssa1 0.61fF
C161 user_analog_project_wrapper_empty_0/gpio_noesd[6] vssa1 0.61fF
C162 user_analog_project_wrapper_empty_0/io_in_3v3[13] vssa1 0.61fF
C163 user_analog_project_wrapper_empty_0/io_in[13] vssa1 0.61fF
C164 user_analog_project_wrapper_empty_0/io_out[13] vssa1 0.61fF
C165 user_analog_project_wrapper_empty_0/io_oeb[13] vssa1 0.61fF
C166 user_analog_project_wrapper_empty_0/vccd1 vssa1 13.04fF
C167 user_analog_project_wrapper_empty_0/vccd2 vssa1 13.04fF
C168 user_analog_project_wrapper_empty_0/io_analog[0] vssa1 6.83fF
C169 user_analog_project_wrapper_empty_0/io_analog[10] vssa1 6.83fF
C170 user_analog_project_wrapper_empty_0/io_clamp_high[0] vssa1 3.58fF
C171 user_analog_project_wrapper_empty_0/io_clamp_low[0] vssa1 3.58fF
C172 user_analog_project_wrapper_empty_0/io_clamp_high[1] vssa1 3.58fF
C173 user_analog_project_wrapper_empty_0/io_clamp_low[1] vssa1 3.58fF
C174 user_analog_project_wrapper_empty_0/io_clamp_high[2] vssa1 3.58fF
C175 user_analog_project_wrapper_empty_0/io_clamp_low[2] vssa1 3.58fF
C176 user_analog_project_wrapper_empty_0/io_analog[7] vssa1 6.83fF
C177 user_analog_project_wrapper_empty_0/io_analog[8] vssa1 6.83fF
C178 user_analog_project_wrapper_empty_0/io_analog[9] vssa1 6.83fF
C179 user_analog_project_wrapper_empty_0/user_irq[2] vssa1 0.63fF
C180 user_analog_project_wrapper_empty_0/user_irq[1] vssa1 0.63fF
C181 user_analog_project_wrapper_empty_0/user_irq[0] vssa1 0.63fF
C182 user_analog_project_wrapper_empty_0/user_clock2 vssa1 0.63fF
C183 user_analog_project_wrapper_empty_0/la_oenb[127] vssa1 0.63fF
C184 user_analog_project_wrapper_empty_0/la_data_out[127] vssa1 0.63fF
C185 user_analog_project_wrapper_empty_0/la_data_in[127] vssa1 0.63fF
C186 user_analog_project_wrapper_empty_0/la_oenb[126] vssa1 0.63fF
C187 user_analog_project_wrapper_empty_0/la_data_out[126] vssa1 0.63fF
C188 user_analog_project_wrapper_empty_0/la_data_in[126] vssa1 0.63fF
C189 user_analog_project_wrapper_empty_0/la_oenb[125] vssa1 0.63fF
C190 user_analog_project_wrapper_empty_0/la_data_out[125] vssa1 0.63fF
C191 user_analog_project_wrapper_empty_0/la_data_in[125] vssa1 0.63fF
C192 user_analog_project_wrapper_empty_0/la_oenb[124] vssa1 0.63fF
C193 user_analog_project_wrapper_empty_0/la_data_out[124] vssa1 0.63fF
C194 user_analog_project_wrapper_empty_0/la_data_in[124] vssa1 0.63fF
C195 user_analog_project_wrapper_empty_0/la_oenb[123] vssa1 0.63fF
C196 user_analog_project_wrapper_empty_0/la_data_out[123] vssa1 0.63fF
C197 user_analog_project_wrapper_empty_0/la_data_in[123] vssa1 0.63fF
C198 user_analog_project_wrapper_empty_0/la_oenb[122] vssa1 0.63fF
C199 user_analog_project_wrapper_empty_0/la_data_out[122] vssa1 0.63fF
C200 user_analog_project_wrapper_empty_0/la_data_in[122] vssa1 0.63fF
C201 user_analog_project_wrapper_empty_0/la_oenb[121] vssa1 0.63fF
C202 user_analog_project_wrapper_empty_0/la_data_out[121] vssa1 0.63fF
C203 user_analog_project_wrapper_empty_0/la_data_in[121] vssa1 0.63fF
C204 user_analog_project_wrapper_empty_0/la_oenb[120] vssa1 0.63fF
C205 user_analog_project_wrapper_empty_0/la_data_out[120] vssa1 0.63fF
C206 user_analog_project_wrapper_empty_0/la_data_in[120] vssa1 0.63fF
C207 user_analog_project_wrapper_empty_0/la_oenb[119] vssa1 0.63fF
C208 user_analog_project_wrapper_empty_0/la_data_out[119] vssa1 0.63fF
C209 user_analog_project_wrapper_empty_0/la_data_in[119] vssa1 0.63fF
C210 user_analog_project_wrapper_empty_0/la_oenb[118] vssa1 0.63fF
C211 user_analog_project_wrapper_empty_0/la_data_out[118] vssa1 0.63fF
C212 user_analog_project_wrapper_empty_0/la_data_in[118] vssa1 0.63fF
C213 user_analog_project_wrapper_empty_0/la_oenb[117] vssa1 0.63fF
C214 user_analog_project_wrapper_empty_0/la_data_out[117] vssa1 0.63fF
C215 user_analog_project_wrapper_empty_0/la_data_in[117] vssa1 0.63fF
C216 user_analog_project_wrapper_empty_0/la_oenb[116] vssa1 0.63fF
C217 user_analog_project_wrapper_empty_0/la_data_out[116] vssa1 0.63fF
C218 user_analog_project_wrapper_empty_0/la_data_in[116] vssa1 0.63fF
C219 user_analog_project_wrapper_empty_0/la_oenb[115] vssa1 0.63fF
C220 user_analog_project_wrapper_empty_0/la_data_out[115] vssa1 0.63fF
C221 user_analog_project_wrapper_empty_0/la_data_in[115] vssa1 0.63fF
C222 user_analog_project_wrapper_empty_0/la_oenb[114] vssa1 0.63fF
C223 user_analog_project_wrapper_empty_0/la_data_out[114] vssa1 0.63fF
C224 user_analog_project_wrapper_empty_0/la_data_in[114] vssa1 0.63fF
C225 user_analog_project_wrapper_empty_0/la_oenb[113] vssa1 0.63fF
C226 user_analog_project_wrapper_empty_0/la_data_out[113] vssa1 0.63fF
C227 user_analog_project_wrapper_empty_0/la_data_in[113] vssa1 0.63fF
C228 user_analog_project_wrapper_empty_0/la_oenb[112] vssa1 0.63fF
C229 user_analog_project_wrapper_empty_0/la_data_out[112] vssa1 0.63fF
C230 user_analog_project_wrapper_empty_0/la_data_in[112] vssa1 0.63fF
C231 user_analog_project_wrapper_empty_0/la_oenb[111] vssa1 0.63fF
C232 user_analog_project_wrapper_empty_0/la_data_out[111] vssa1 0.63fF
C233 user_analog_project_wrapper_empty_0/la_data_in[111] vssa1 0.63fF
C234 user_analog_project_wrapper_empty_0/la_oenb[110] vssa1 0.63fF
C235 user_analog_project_wrapper_empty_0/la_data_out[110] vssa1 0.63fF
C236 user_analog_project_wrapper_empty_0/la_data_in[110] vssa1 0.63fF
C237 user_analog_project_wrapper_empty_0/la_oenb[109] vssa1 0.63fF
C238 user_analog_project_wrapper_empty_0/la_data_out[109] vssa1 0.63fF
C239 user_analog_project_wrapper_empty_0/la_data_in[109] vssa1 0.63fF
C240 user_analog_project_wrapper_empty_0/la_oenb[108] vssa1 0.63fF
C241 user_analog_project_wrapper_empty_0/la_data_out[108] vssa1 0.63fF
C242 user_analog_project_wrapper_empty_0/la_data_in[108] vssa1 0.63fF
C243 user_analog_project_wrapper_empty_0/la_oenb[107] vssa1 0.63fF
C244 user_analog_project_wrapper_empty_0/la_data_out[107] vssa1 0.63fF
C245 user_analog_project_wrapper_empty_0/la_data_in[107] vssa1 0.63fF
C246 user_analog_project_wrapper_empty_0/la_oenb[106] vssa1 0.63fF
C247 user_analog_project_wrapper_empty_0/la_data_out[106] vssa1 0.63fF
C248 user_analog_project_wrapper_empty_0/la_data_in[106] vssa1 0.63fF
C249 user_analog_project_wrapper_empty_0/la_oenb[105] vssa1 0.63fF
C250 user_analog_project_wrapper_empty_0/la_data_out[105] vssa1 0.63fF
C251 user_analog_project_wrapper_empty_0/la_data_in[105] vssa1 0.63fF
C252 user_analog_project_wrapper_empty_0/la_oenb[104] vssa1 0.63fF
C253 user_analog_project_wrapper_empty_0/la_data_out[104] vssa1 0.63fF
C254 user_analog_project_wrapper_empty_0/la_data_in[104] vssa1 0.63fF
C255 user_analog_project_wrapper_empty_0/la_oenb[103] vssa1 0.63fF
C256 user_analog_project_wrapper_empty_0/la_data_out[103] vssa1 0.63fF
C257 user_analog_project_wrapper_empty_0/la_data_in[103] vssa1 0.63fF
C258 user_analog_project_wrapper_empty_0/la_oenb[102] vssa1 0.63fF
C259 user_analog_project_wrapper_empty_0/la_data_out[102] vssa1 0.63fF
C260 user_analog_project_wrapper_empty_0/la_data_in[102] vssa1 0.63fF
C261 user_analog_project_wrapper_empty_0/la_oenb[101] vssa1 0.63fF
C262 user_analog_project_wrapper_empty_0/la_data_out[101] vssa1 0.63fF
C263 user_analog_project_wrapper_empty_0/la_data_in[101] vssa1 0.63fF
C264 user_analog_project_wrapper_empty_0/la_oenb[100] vssa1 0.63fF
C265 user_analog_project_wrapper_empty_0/la_data_out[100] vssa1 0.63fF
C266 user_analog_project_wrapper_empty_0/la_data_in[100] vssa1 0.63fF
C267 user_analog_project_wrapper_empty_0/la_oenb[99] vssa1 0.63fF
C268 user_analog_project_wrapper_empty_0/la_data_out[99] vssa1 0.63fF
C269 user_analog_project_wrapper_empty_0/la_data_in[99] vssa1 0.63fF
C270 user_analog_project_wrapper_empty_0/la_oenb[98] vssa1 0.63fF
C271 user_analog_project_wrapper_empty_0/la_data_out[98] vssa1 0.63fF
C272 user_analog_project_wrapper_empty_0/la_data_in[98] vssa1 0.63fF
C273 user_analog_project_wrapper_empty_0/la_oenb[97] vssa1 0.63fF
C274 user_analog_project_wrapper_empty_0/la_data_out[97] vssa1 0.63fF
C275 user_analog_project_wrapper_empty_0/la_data_in[97] vssa1 0.63fF
C276 user_analog_project_wrapper_empty_0/la_oenb[96] vssa1 0.63fF
C277 user_analog_project_wrapper_empty_0/la_data_out[96] vssa1 0.63fF
C278 user_analog_project_wrapper_empty_0/la_data_in[96] vssa1 0.63fF
C279 user_analog_project_wrapper_empty_0/la_oenb[95] vssa1 0.63fF
C280 user_analog_project_wrapper_empty_0/la_data_out[95] vssa1 0.63fF
C281 user_analog_project_wrapper_empty_0/la_data_in[95] vssa1 0.63fF
C282 user_analog_project_wrapper_empty_0/la_oenb[94] vssa1 0.63fF
C283 user_analog_project_wrapper_empty_0/la_data_out[94] vssa1 0.63fF
C284 user_analog_project_wrapper_empty_0/la_data_in[94] vssa1 0.63fF
C285 user_analog_project_wrapper_empty_0/la_oenb[93] vssa1 0.63fF
C286 user_analog_project_wrapper_empty_0/la_data_out[93] vssa1 0.63fF
C287 user_analog_project_wrapper_empty_0/la_data_in[93] vssa1 0.63fF
C288 user_analog_project_wrapper_empty_0/la_oenb[92] vssa1 0.63fF
C289 user_analog_project_wrapper_empty_0/la_data_out[92] vssa1 0.63fF
C290 user_analog_project_wrapper_empty_0/la_data_in[92] vssa1 0.63fF
C291 user_analog_project_wrapper_empty_0/la_oenb[91] vssa1 0.63fF
C292 user_analog_project_wrapper_empty_0/la_data_out[91] vssa1 0.63fF
C293 user_analog_project_wrapper_empty_0/la_data_in[91] vssa1 0.63fF
C294 user_analog_project_wrapper_empty_0/la_oenb[90] vssa1 0.63fF
C295 user_analog_project_wrapper_empty_0/la_data_out[90] vssa1 0.63fF
C296 user_analog_project_wrapper_empty_0/la_data_in[90] vssa1 0.63fF
C297 user_analog_project_wrapper_empty_0/la_oenb[89] vssa1 0.63fF
C298 user_analog_project_wrapper_empty_0/la_data_out[89] vssa1 0.63fF
C299 user_analog_project_wrapper_empty_0/la_data_in[89] vssa1 0.63fF
C300 user_analog_project_wrapper_empty_0/la_oenb[88] vssa1 0.63fF
C301 user_analog_project_wrapper_empty_0/la_data_out[88] vssa1 0.63fF
C302 user_analog_project_wrapper_empty_0/la_data_in[88] vssa1 0.63fF
C303 user_analog_project_wrapper_empty_0/la_oenb[87] vssa1 0.63fF
C304 user_analog_project_wrapper_empty_0/la_data_out[87] vssa1 0.63fF
C305 user_analog_project_wrapper_empty_0/la_data_in[87] vssa1 0.63fF
C306 user_analog_project_wrapper_empty_0/la_oenb[86] vssa1 0.63fF
C307 user_analog_project_wrapper_empty_0/la_data_out[86] vssa1 0.63fF
C308 user_analog_project_wrapper_empty_0/la_data_in[86] vssa1 0.63fF
C309 user_analog_project_wrapper_empty_0/la_oenb[85] vssa1 0.63fF
C310 user_analog_project_wrapper_empty_0/la_data_out[85] vssa1 0.63fF
C311 user_analog_project_wrapper_empty_0/la_data_in[85] vssa1 0.63fF
C312 user_analog_project_wrapper_empty_0/la_oenb[84] vssa1 0.63fF
C313 user_analog_project_wrapper_empty_0/la_data_out[84] vssa1 0.63fF
C314 user_analog_project_wrapper_empty_0/la_data_in[84] vssa1 0.63fF
C315 user_analog_project_wrapper_empty_0/la_oenb[83] vssa1 0.63fF
C316 user_analog_project_wrapper_empty_0/la_data_out[83] vssa1 0.63fF
C317 user_analog_project_wrapper_empty_0/la_data_in[83] vssa1 0.63fF
C318 user_analog_project_wrapper_empty_0/la_oenb[82] vssa1 0.63fF
C319 user_analog_project_wrapper_empty_0/la_data_out[82] vssa1 0.63fF
C320 user_analog_project_wrapper_empty_0/la_data_in[82] vssa1 0.63fF
C321 user_analog_project_wrapper_empty_0/la_oenb[81] vssa1 0.63fF
C322 user_analog_project_wrapper_empty_0/la_data_out[81] vssa1 0.63fF
C323 user_analog_project_wrapper_empty_0/la_data_in[81] vssa1 0.63fF
C324 user_analog_project_wrapper_empty_0/la_oenb[80] vssa1 0.63fF
C325 user_analog_project_wrapper_empty_0/la_data_out[80] vssa1 0.63fF
C326 user_analog_project_wrapper_empty_0/la_data_in[80] vssa1 0.63fF
C327 user_analog_project_wrapper_empty_0/la_oenb[79] vssa1 0.63fF
C328 user_analog_project_wrapper_empty_0/la_data_out[79] vssa1 0.63fF
C329 user_analog_project_wrapper_empty_0/la_data_in[79] vssa1 0.63fF
C330 user_analog_project_wrapper_empty_0/la_oenb[78] vssa1 0.63fF
C331 user_analog_project_wrapper_empty_0/la_data_out[78] vssa1 0.63fF
C332 user_analog_project_wrapper_empty_0/la_data_in[78] vssa1 0.63fF
C333 user_analog_project_wrapper_empty_0/la_oenb[77] vssa1 0.63fF
C334 user_analog_project_wrapper_empty_0/la_data_out[77] vssa1 0.63fF
C335 user_analog_project_wrapper_empty_0/la_data_in[77] vssa1 0.63fF
C336 user_analog_project_wrapper_empty_0/la_oenb[76] vssa1 0.63fF
C337 user_analog_project_wrapper_empty_0/la_data_out[76] vssa1 0.63fF
C338 user_analog_project_wrapper_empty_0/la_data_in[76] vssa1 0.63fF
C339 user_analog_project_wrapper_empty_0/la_oenb[75] vssa1 0.63fF
C340 user_analog_project_wrapper_empty_0/la_data_out[75] vssa1 0.63fF
C341 user_analog_project_wrapper_empty_0/la_data_in[75] vssa1 0.63fF
C342 user_analog_project_wrapper_empty_0/la_oenb[74] vssa1 0.63fF
C343 user_analog_project_wrapper_empty_0/la_data_out[74] vssa1 0.63fF
C344 user_analog_project_wrapper_empty_0/la_data_in[74] vssa1 0.63fF
C345 user_analog_project_wrapper_empty_0/la_oenb[73] vssa1 0.63fF
C346 user_analog_project_wrapper_empty_0/la_data_out[73] vssa1 0.63fF
C347 user_analog_project_wrapper_empty_0/la_data_in[73] vssa1 0.63fF
C348 user_analog_project_wrapper_empty_0/la_oenb[72] vssa1 0.63fF
C349 user_analog_project_wrapper_empty_0/la_data_out[72] vssa1 0.63fF
C350 user_analog_project_wrapper_empty_0/la_data_in[72] vssa1 0.63fF
C351 user_analog_project_wrapper_empty_0/la_oenb[71] vssa1 0.63fF
C352 user_analog_project_wrapper_empty_0/la_data_out[71] vssa1 0.63fF
C353 user_analog_project_wrapper_empty_0/la_data_in[71] vssa1 0.63fF
C354 user_analog_project_wrapper_empty_0/la_oenb[70] vssa1 0.63fF
C355 user_analog_project_wrapper_empty_0/la_data_out[70] vssa1 0.63fF
C356 user_analog_project_wrapper_empty_0/la_data_in[70] vssa1 0.63fF
C357 user_analog_project_wrapper_empty_0/la_oenb[69] vssa1 0.63fF
C358 user_analog_project_wrapper_empty_0/la_data_out[69] vssa1 0.63fF
C359 user_analog_project_wrapper_empty_0/la_data_in[69] vssa1 0.63fF
C360 user_analog_project_wrapper_empty_0/la_oenb[68] vssa1 0.63fF
C361 user_analog_project_wrapper_empty_0/la_data_out[68] vssa1 0.63fF
C362 user_analog_project_wrapper_empty_0/la_data_in[68] vssa1 0.63fF
C363 user_analog_project_wrapper_empty_0/la_oenb[67] vssa1 0.63fF
C364 user_analog_project_wrapper_empty_0/la_data_out[67] vssa1 0.63fF
C365 user_analog_project_wrapper_empty_0/la_data_in[67] vssa1 0.63fF
C366 user_analog_project_wrapper_empty_0/la_oenb[66] vssa1 0.63fF
C367 user_analog_project_wrapper_empty_0/la_data_out[66] vssa1 0.63fF
C368 user_analog_project_wrapper_empty_0/la_data_in[66] vssa1 0.63fF
C369 user_analog_project_wrapper_empty_0/la_oenb[65] vssa1 0.63fF
C370 user_analog_project_wrapper_empty_0/la_data_out[65] vssa1 0.63fF
C371 user_analog_project_wrapper_empty_0/la_data_in[65] vssa1 0.63fF
C372 user_analog_project_wrapper_empty_0/la_oenb[64] vssa1 0.63fF
C373 user_analog_project_wrapper_empty_0/la_data_out[64] vssa1 0.63fF
C374 user_analog_project_wrapper_empty_0/la_data_in[64] vssa1 0.63fF
C375 user_analog_project_wrapper_empty_0/la_oenb[63] vssa1 0.63fF
C376 user_analog_project_wrapper_empty_0/la_data_out[63] vssa1 0.63fF
C377 user_analog_project_wrapper_empty_0/la_data_in[63] vssa1 0.63fF
C378 user_analog_project_wrapper_empty_0/la_oenb[62] vssa1 0.63fF
C379 user_analog_project_wrapper_empty_0/la_data_out[62] vssa1 0.63fF
C380 user_analog_project_wrapper_empty_0/la_data_in[62] vssa1 0.63fF
C381 user_analog_project_wrapper_empty_0/la_oenb[61] vssa1 0.63fF
C382 user_analog_project_wrapper_empty_0/la_data_out[61] vssa1 0.63fF
C383 user_analog_project_wrapper_empty_0/la_data_in[61] vssa1 0.63fF
C384 user_analog_project_wrapper_empty_0/la_oenb[60] vssa1 0.63fF
C385 user_analog_project_wrapper_empty_0/la_data_out[60] vssa1 0.63fF
C386 user_analog_project_wrapper_empty_0/la_data_in[60] vssa1 0.63fF
C387 user_analog_project_wrapper_empty_0/la_oenb[59] vssa1 0.63fF
C388 user_analog_project_wrapper_empty_0/la_data_out[59] vssa1 0.63fF
C389 user_analog_project_wrapper_empty_0/la_data_in[59] vssa1 0.63fF
C390 user_analog_project_wrapper_empty_0/la_oenb[58] vssa1 0.63fF
C391 user_analog_project_wrapper_empty_0/la_data_out[58] vssa1 0.63fF
C392 user_analog_project_wrapper_empty_0/la_data_in[58] vssa1 0.63fF
C393 user_analog_project_wrapper_empty_0/la_oenb[57] vssa1 0.63fF
C394 user_analog_project_wrapper_empty_0/la_data_out[57] vssa1 0.63fF
C395 user_analog_project_wrapper_empty_0/la_data_in[57] vssa1 0.63fF
C396 user_analog_project_wrapper_empty_0/la_oenb[56] vssa1 0.63fF
C397 user_analog_project_wrapper_empty_0/la_data_out[56] vssa1 0.63fF
C398 user_analog_project_wrapper_empty_0/la_data_in[56] vssa1 0.63fF
C399 user_analog_project_wrapper_empty_0/la_oenb[55] vssa1 0.63fF
C400 user_analog_project_wrapper_empty_0/la_data_out[55] vssa1 0.63fF
C401 user_analog_project_wrapper_empty_0/la_data_in[55] vssa1 0.63fF
C402 user_analog_project_wrapper_empty_0/la_oenb[54] vssa1 0.63fF
C403 user_analog_project_wrapper_empty_0/la_data_out[54] vssa1 0.63fF
C404 user_analog_project_wrapper_empty_0/la_data_in[54] vssa1 0.63fF
C405 user_analog_project_wrapper_empty_0/la_oenb[53] vssa1 0.63fF
C406 user_analog_project_wrapper_empty_0/la_data_out[53] vssa1 0.63fF
C407 user_analog_project_wrapper_empty_0/la_data_in[53] vssa1 0.63fF
C408 user_analog_project_wrapper_empty_0/la_oenb[52] vssa1 0.63fF
C409 user_analog_project_wrapper_empty_0/la_data_out[52] vssa1 0.63fF
C410 user_analog_project_wrapper_empty_0/la_data_in[52] vssa1 0.63fF
C411 user_analog_project_wrapper_empty_0/la_oenb[51] vssa1 0.63fF
C412 user_analog_project_wrapper_empty_0/la_data_out[51] vssa1 0.63fF
C413 user_analog_project_wrapper_empty_0/la_data_in[51] vssa1 0.63fF
C414 user_analog_project_wrapper_empty_0/la_oenb[50] vssa1 0.63fF
C415 user_analog_project_wrapper_empty_0/la_data_out[50] vssa1 0.63fF
C416 user_analog_project_wrapper_empty_0/la_data_in[50] vssa1 0.63fF
C417 user_analog_project_wrapper_empty_0/la_oenb[49] vssa1 0.63fF
C418 user_analog_project_wrapper_empty_0/la_data_out[49] vssa1 0.63fF
C419 user_analog_project_wrapper_empty_0/la_data_in[49] vssa1 0.63fF
C420 user_analog_project_wrapper_empty_0/la_oenb[48] vssa1 0.63fF
C421 user_analog_project_wrapper_empty_0/la_data_out[48] vssa1 0.63fF
C422 user_analog_project_wrapper_empty_0/la_data_in[48] vssa1 0.63fF
C423 user_analog_project_wrapper_empty_0/la_oenb[47] vssa1 0.63fF
C424 user_analog_project_wrapper_empty_0/la_data_out[47] vssa1 0.63fF
C425 user_analog_project_wrapper_empty_0/la_data_in[47] vssa1 0.63fF
C426 user_analog_project_wrapper_empty_0/la_oenb[46] vssa1 0.63fF
C427 user_analog_project_wrapper_empty_0/la_data_out[46] vssa1 0.63fF
C428 user_analog_project_wrapper_empty_0/la_data_in[46] vssa1 0.63fF
C429 user_analog_project_wrapper_empty_0/la_oenb[45] vssa1 0.63fF
C430 user_analog_project_wrapper_empty_0/la_data_out[45] vssa1 0.63fF
C431 user_analog_project_wrapper_empty_0/la_data_in[45] vssa1 0.63fF
C432 user_analog_project_wrapper_empty_0/la_oenb[44] vssa1 0.63fF
C433 user_analog_project_wrapper_empty_0/la_data_out[44] vssa1 0.63fF
C434 user_analog_project_wrapper_empty_0/la_data_in[44] vssa1 0.63fF
C435 user_analog_project_wrapper_empty_0/la_oenb[43] vssa1 0.63fF
C436 user_analog_project_wrapper_empty_0/la_data_out[43] vssa1 0.63fF
C437 user_analog_project_wrapper_empty_0/la_data_in[43] vssa1 0.63fF
C438 user_analog_project_wrapper_empty_0/la_oenb[42] vssa1 0.63fF
C439 user_analog_project_wrapper_empty_0/la_data_out[42] vssa1 0.63fF
C440 user_analog_project_wrapper_empty_0/la_data_in[42] vssa1 0.63fF
C441 user_analog_project_wrapper_empty_0/la_oenb[41] vssa1 0.63fF
C442 user_analog_project_wrapper_empty_0/la_data_out[41] vssa1 0.63fF
C443 user_analog_project_wrapper_empty_0/la_data_in[41] vssa1 0.63fF
C444 user_analog_project_wrapper_empty_0/la_oenb[40] vssa1 0.63fF
C445 user_analog_project_wrapper_empty_0/la_data_out[40] vssa1 0.63fF
C446 user_analog_project_wrapper_empty_0/la_data_in[40] vssa1 0.63fF
C447 user_analog_project_wrapper_empty_0/la_oenb[39] vssa1 0.63fF
C448 user_analog_project_wrapper_empty_0/la_data_out[39] vssa1 0.63fF
C449 user_analog_project_wrapper_empty_0/la_data_in[39] vssa1 0.63fF
C450 user_analog_project_wrapper_empty_0/la_oenb[38] vssa1 0.63fF
C451 user_analog_project_wrapper_empty_0/la_data_out[38] vssa1 0.63fF
C452 user_analog_project_wrapper_empty_0/la_data_in[38] vssa1 0.63fF
C453 user_analog_project_wrapper_empty_0/la_oenb[37] vssa1 0.63fF
C454 user_analog_project_wrapper_empty_0/la_data_out[37] vssa1 0.63fF
C455 user_analog_project_wrapper_empty_0/la_data_in[37] vssa1 0.63fF
C456 user_analog_project_wrapper_empty_0/la_oenb[36] vssa1 0.63fF
C457 user_analog_project_wrapper_empty_0/la_data_out[36] vssa1 0.63fF
C458 user_analog_project_wrapper_empty_0/la_data_in[36] vssa1 0.63fF
C459 user_analog_project_wrapper_empty_0/la_oenb[35] vssa1 0.63fF
C460 user_analog_project_wrapper_empty_0/la_data_out[35] vssa1 0.63fF
C461 user_analog_project_wrapper_empty_0/la_data_in[35] vssa1 0.63fF
C462 user_analog_project_wrapper_empty_0/la_oenb[34] vssa1 0.63fF
C463 user_analog_project_wrapper_empty_0/la_data_out[34] vssa1 0.63fF
C464 user_analog_project_wrapper_empty_0/la_data_in[34] vssa1 0.63fF
C465 user_analog_project_wrapper_empty_0/la_oenb[33] vssa1 0.63fF
C466 user_analog_project_wrapper_empty_0/la_data_out[33] vssa1 0.63fF
C467 user_analog_project_wrapper_empty_0/la_data_in[33] vssa1 0.63fF
C468 user_analog_project_wrapper_empty_0/la_oenb[32] vssa1 0.63fF
C469 user_analog_project_wrapper_empty_0/la_data_out[32] vssa1 0.63fF
C470 user_analog_project_wrapper_empty_0/la_data_in[32] vssa1 0.63fF
C471 user_analog_project_wrapper_empty_0/la_oenb[31] vssa1 0.63fF
C472 user_analog_project_wrapper_empty_0/la_data_out[31] vssa1 0.63fF
C473 user_analog_project_wrapper_empty_0/la_data_in[31] vssa1 0.63fF
C474 user_analog_project_wrapper_empty_0/la_oenb[30] vssa1 0.63fF
C475 user_analog_project_wrapper_empty_0/la_data_out[30] vssa1 0.63fF
C476 user_analog_project_wrapper_empty_0/la_data_in[30] vssa1 0.63fF
C477 user_analog_project_wrapper_empty_0/la_oenb[29] vssa1 0.63fF
C478 user_analog_project_wrapper_empty_0/la_data_out[29] vssa1 0.63fF
C479 user_analog_project_wrapper_empty_0/la_data_in[29] vssa1 0.63fF
C480 user_analog_project_wrapper_empty_0/la_oenb[28] vssa1 0.63fF
C481 user_analog_project_wrapper_empty_0/la_data_out[28] vssa1 0.63fF
C482 user_analog_project_wrapper_empty_0/la_data_in[28] vssa1 0.63fF
C483 user_analog_project_wrapper_empty_0/la_oenb[27] vssa1 0.63fF
C484 user_analog_project_wrapper_empty_0/la_data_out[27] vssa1 0.63fF
C485 user_analog_project_wrapper_empty_0/la_data_in[27] vssa1 0.63fF
C486 user_analog_project_wrapper_empty_0/la_oenb[26] vssa1 0.63fF
C487 user_analog_project_wrapper_empty_0/la_data_out[26] vssa1 0.63fF
C488 user_analog_project_wrapper_empty_0/la_data_in[26] vssa1 0.63fF
C489 user_analog_project_wrapper_empty_0/la_oenb[25] vssa1 0.63fF
C490 user_analog_project_wrapper_empty_0/la_data_out[25] vssa1 0.63fF
C491 user_analog_project_wrapper_empty_0/la_data_in[25] vssa1 0.63fF
C492 user_analog_project_wrapper_empty_0/la_oenb[24] vssa1 0.63fF
C493 user_analog_project_wrapper_empty_0/la_data_out[24] vssa1 0.63fF
C494 user_analog_project_wrapper_empty_0/la_data_in[24] vssa1 0.63fF
C495 user_analog_project_wrapper_empty_0/la_oenb[23] vssa1 0.63fF
C496 user_analog_project_wrapper_empty_0/la_data_out[23] vssa1 0.63fF
C497 user_analog_project_wrapper_empty_0/la_data_in[23] vssa1 0.63fF
C498 user_analog_project_wrapper_empty_0/la_oenb[22] vssa1 0.63fF
C499 user_analog_project_wrapper_empty_0/la_data_out[22] vssa1 0.63fF
C500 user_analog_project_wrapper_empty_0/la_data_in[22] vssa1 0.63fF
C501 user_analog_project_wrapper_empty_0/la_oenb[21] vssa1 0.63fF
C502 user_analog_project_wrapper_empty_0/la_data_out[21] vssa1 0.63fF
C503 user_analog_project_wrapper_empty_0/la_data_in[21] vssa1 0.63fF
C504 user_analog_project_wrapper_empty_0/la_oenb[20] vssa1 0.63fF
C505 user_analog_project_wrapper_empty_0/la_data_out[20] vssa1 0.63fF
C506 user_analog_project_wrapper_empty_0/la_data_in[20] vssa1 0.63fF
C507 user_analog_project_wrapper_empty_0/la_oenb[19] vssa1 0.63fF
C508 user_analog_project_wrapper_empty_0/la_data_out[19] vssa1 0.63fF
C509 user_analog_project_wrapper_empty_0/la_data_in[19] vssa1 0.63fF
C510 user_analog_project_wrapper_empty_0/la_oenb[18] vssa1 0.63fF
C511 user_analog_project_wrapper_empty_0/la_data_out[18] vssa1 0.63fF
C512 user_analog_project_wrapper_empty_0/la_data_in[18] vssa1 0.63fF
C513 user_analog_project_wrapper_empty_0/la_oenb[17] vssa1 0.63fF
C514 user_analog_project_wrapper_empty_0/la_data_out[17] vssa1 0.63fF
C515 user_analog_project_wrapper_empty_0/la_data_in[17] vssa1 0.63fF
C516 user_analog_project_wrapper_empty_0/la_oenb[16] vssa1 0.63fF
C517 user_analog_project_wrapper_empty_0/la_data_out[16] vssa1 0.63fF
C518 user_analog_project_wrapper_empty_0/la_data_in[16] vssa1 0.63fF
C519 user_analog_project_wrapper_empty_0/la_oenb[15] vssa1 0.63fF
C520 user_analog_project_wrapper_empty_0/la_data_out[15] vssa1 0.63fF
C521 user_analog_project_wrapper_empty_0/la_data_in[15] vssa1 0.63fF
C522 user_analog_project_wrapper_empty_0/la_oenb[14] vssa1 0.63fF
C523 user_analog_project_wrapper_empty_0/la_data_out[14] vssa1 0.63fF
C524 user_analog_project_wrapper_empty_0/la_data_in[14] vssa1 0.63fF
C525 user_analog_project_wrapper_empty_0/la_oenb[13] vssa1 0.63fF
C526 user_analog_project_wrapper_empty_0/la_data_out[13] vssa1 0.63fF
C527 user_analog_project_wrapper_empty_0/la_data_in[13] vssa1 0.63fF
C528 user_analog_project_wrapper_empty_0/la_oenb[12] vssa1 0.63fF
C529 user_analog_project_wrapper_empty_0/la_data_out[12] vssa1 0.63fF
C530 user_analog_project_wrapper_empty_0/la_data_in[12] vssa1 0.63fF
C531 user_analog_project_wrapper_empty_0/la_oenb[11] vssa1 0.63fF
C532 user_analog_project_wrapper_empty_0/la_data_out[11] vssa1 0.63fF
C533 user_analog_project_wrapper_empty_0/la_data_in[11] vssa1 0.63fF
C534 user_analog_project_wrapper_empty_0/la_oenb[10] vssa1 0.63fF
C535 user_analog_project_wrapper_empty_0/la_data_out[10] vssa1 0.63fF
C536 user_analog_project_wrapper_empty_0/la_data_in[10] vssa1 0.63fF
C537 user_analog_project_wrapper_empty_0/la_oenb[9] vssa1 0.63fF
C538 user_analog_project_wrapper_empty_0/la_data_out[9] vssa1 0.63fF
C539 user_analog_project_wrapper_empty_0/la_data_in[9] vssa1 0.63fF
C540 user_analog_project_wrapper_empty_0/la_oenb[8] vssa1 0.63fF
C541 user_analog_project_wrapper_empty_0/la_data_out[8] vssa1 0.63fF
C542 user_analog_project_wrapper_empty_0/la_data_in[8] vssa1 0.63fF
C543 user_analog_project_wrapper_empty_0/la_oenb[7] vssa1 0.63fF
C544 user_analog_project_wrapper_empty_0/la_data_out[7] vssa1 0.63fF
C545 user_analog_project_wrapper_empty_0/la_data_in[7] vssa1 0.63fF
C546 user_analog_project_wrapper_empty_0/la_oenb[6] vssa1 0.63fF
C547 user_analog_project_wrapper_empty_0/la_data_out[6] vssa1 0.63fF
C548 user_analog_project_wrapper_empty_0/la_data_in[6] vssa1 0.63fF
C549 user_analog_project_wrapper_empty_0/la_oenb[5] vssa1 0.63fF
C550 user_analog_project_wrapper_empty_0/la_data_out[5] vssa1 0.63fF
C551 user_analog_project_wrapper_empty_0/la_data_in[5] vssa1 0.63fF
C552 user_analog_project_wrapper_empty_0/la_oenb[4] vssa1 0.63fF
C553 user_analog_project_wrapper_empty_0/la_data_out[4] vssa1 0.63fF
C554 user_analog_project_wrapper_empty_0/la_data_in[4] vssa1 0.63fF
C555 user_analog_project_wrapper_empty_0/la_oenb[3] vssa1 0.63fF
C556 user_analog_project_wrapper_empty_0/la_data_out[3] vssa1 0.63fF
C557 user_analog_project_wrapper_empty_0/la_data_in[3] vssa1 0.63fF
C558 user_analog_project_wrapper_empty_0/la_oenb[2] vssa1 0.63fF
C559 user_analog_project_wrapper_empty_0/la_data_out[2] vssa1 0.63fF
C560 user_analog_project_wrapper_empty_0/la_data_in[2] vssa1 0.63fF
C561 user_analog_project_wrapper_empty_0/la_oenb[1] vssa1 0.63fF
C562 user_analog_project_wrapper_empty_0/la_data_out[1] vssa1 0.63fF
C563 user_analog_project_wrapper_empty_0/la_data_in[1] vssa1 0.63fF
C564 user_analog_project_wrapper_empty_0/la_oenb[0] vssa1 0.63fF
C565 user_analog_project_wrapper_empty_0/la_data_out[0] vssa1 0.63fF
C566 user_analog_project_wrapper_empty_0/la_data_in[0] vssa1 0.63fF
C567 user_analog_project_wrapper_empty_0/wbs_dat_o[31] vssa1 0.63fF
C568 user_analog_project_wrapper_empty_0/wbs_dat_i[31] vssa1 0.63fF
C569 user_analog_project_wrapper_empty_0/wbs_adr_i[31] vssa1 0.63fF
C570 user_analog_project_wrapper_empty_0/wbs_dat_o[30] vssa1 0.63fF
C571 user_analog_project_wrapper_empty_0/wbs_dat_i[30] vssa1 0.63fF
C572 user_analog_project_wrapper_empty_0/wbs_adr_i[30] vssa1 0.63fF
C573 user_analog_project_wrapper_empty_0/wbs_dat_o[29] vssa1 0.63fF
C574 user_analog_project_wrapper_empty_0/wbs_dat_i[29] vssa1 0.63fF
C575 user_analog_project_wrapper_empty_0/wbs_adr_i[29] vssa1 0.63fF
C576 user_analog_project_wrapper_empty_0/wbs_dat_o[28] vssa1 0.63fF
C577 user_analog_project_wrapper_empty_0/wbs_dat_i[28] vssa1 0.63fF
C578 user_analog_project_wrapper_empty_0/wbs_adr_i[28] vssa1 0.63fF
C579 user_analog_project_wrapper_empty_0/wbs_dat_o[27] vssa1 0.63fF
C580 user_analog_project_wrapper_empty_0/wbs_dat_i[27] vssa1 0.63fF
C581 user_analog_project_wrapper_empty_0/wbs_adr_i[27] vssa1 0.63fF
C582 user_analog_project_wrapper_empty_0/wbs_dat_o[26] vssa1 0.63fF
C583 user_analog_project_wrapper_empty_0/wbs_dat_i[26] vssa1 0.63fF
C584 user_analog_project_wrapper_empty_0/wbs_adr_i[26] vssa1 0.63fF
C585 user_analog_project_wrapper_empty_0/wbs_dat_o[25] vssa1 0.63fF
C586 user_analog_project_wrapper_empty_0/wbs_dat_i[25] vssa1 0.63fF
C587 user_analog_project_wrapper_empty_0/wbs_adr_i[25] vssa1 0.63fF
C588 user_analog_project_wrapper_empty_0/wbs_dat_o[24] vssa1 0.63fF
C589 user_analog_project_wrapper_empty_0/wbs_dat_i[24] vssa1 0.63fF
C590 user_analog_project_wrapper_empty_0/wbs_adr_i[24] vssa1 0.63fF
C591 user_analog_project_wrapper_empty_0/wbs_dat_o[23] vssa1 0.63fF
C592 user_analog_project_wrapper_empty_0/wbs_dat_i[23] vssa1 0.63fF
C593 user_analog_project_wrapper_empty_0/wbs_adr_i[23] vssa1 0.63fF
C594 user_analog_project_wrapper_empty_0/wbs_dat_o[22] vssa1 0.63fF
C595 user_analog_project_wrapper_empty_0/wbs_dat_i[22] vssa1 0.63fF
C596 user_analog_project_wrapper_empty_0/wbs_adr_i[22] vssa1 0.63fF
C597 user_analog_project_wrapper_empty_0/wbs_dat_o[21] vssa1 0.63fF
C598 user_analog_project_wrapper_empty_0/wbs_dat_i[21] vssa1 0.63fF
C599 user_analog_project_wrapper_empty_0/wbs_adr_i[21] vssa1 0.63fF
C600 user_analog_project_wrapper_empty_0/wbs_dat_o[20] vssa1 0.63fF
C601 user_analog_project_wrapper_empty_0/wbs_dat_i[20] vssa1 0.63fF
C602 user_analog_project_wrapper_empty_0/wbs_adr_i[20] vssa1 0.63fF
C603 user_analog_project_wrapper_empty_0/wbs_dat_o[19] vssa1 0.63fF
C604 user_analog_project_wrapper_empty_0/wbs_dat_i[19] vssa1 0.63fF
C605 user_analog_project_wrapper_empty_0/wbs_adr_i[19] vssa1 0.63fF
C606 user_analog_project_wrapper_empty_0/wbs_dat_o[18] vssa1 0.63fF
C607 user_analog_project_wrapper_empty_0/wbs_dat_i[18] vssa1 0.63fF
C608 user_analog_project_wrapper_empty_0/wbs_adr_i[18] vssa1 0.63fF
C609 user_analog_project_wrapper_empty_0/wbs_dat_o[17] vssa1 0.63fF
C610 user_analog_project_wrapper_empty_0/wbs_dat_i[17] vssa1 0.63fF
C611 user_analog_project_wrapper_empty_0/wbs_adr_i[17] vssa1 0.63fF
C612 user_analog_project_wrapper_empty_0/wbs_dat_o[16] vssa1 0.63fF
C613 user_analog_project_wrapper_empty_0/wbs_dat_i[16] vssa1 0.63fF
C614 user_analog_project_wrapper_empty_0/wbs_adr_i[16] vssa1 0.63fF
C615 user_analog_project_wrapper_empty_0/wbs_dat_o[15] vssa1 0.63fF
C616 user_analog_project_wrapper_empty_0/wbs_dat_i[15] vssa1 0.63fF
C617 user_analog_project_wrapper_empty_0/wbs_adr_i[15] vssa1 0.63fF
C618 user_analog_project_wrapper_empty_0/wbs_dat_o[14] vssa1 0.63fF
C619 user_analog_project_wrapper_empty_0/wbs_dat_i[14] vssa1 0.63fF
C620 user_analog_project_wrapper_empty_0/wbs_adr_i[14] vssa1 0.63fF
C621 user_analog_project_wrapper_empty_0/wbs_dat_o[13] vssa1 0.63fF
C622 user_analog_project_wrapper_empty_0/wbs_dat_i[13] vssa1 0.63fF
C623 user_analog_project_wrapper_empty_0/wbs_adr_i[13] vssa1 0.63fF
C624 user_analog_project_wrapper_empty_0/wbs_dat_o[12] vssa1 0.63fF
C625 user_analog_project_wrapper_empty_0/wbs_dat_i[12] vssa1 0.63fF
C626 user_analog_project_wrapper_empty_0/wbs_adr_i[12] vssa1 0.63fF
C627 user_analog_project_wrapper_empty_0/wbs_dat_o[11] vssa1 0.63fF
C628 user_analog_project_wrapper_empty_0/wbs_dat_i[11] vssa1 0.63fF
C629 user_analog_project_wrapper_empty_0/wbs_adr_i[11] vssa1 0.63fF
C630 user_analog_project_wrapper_empty_0/wbs_dat_o[10] vssa1 0.63fF
C631 user_analog_project_wrapper_empty_0/wbs_dat_i[10] vssa1 0.63fF
C632 user_analog_project_wrapper_empty_0/wbs_adr_i[10] vssa1 0.63fF
C633 user_analog_project_wrapper_empty_0/wbs_dat_o[9] vssa1 0.63fF
C634 user_analog_project_wrapper_empty_0/wbs_dat_i[9] vssa1 0.63fF
C635 user_analog_project_wrapper_empty_0/wbs_adr_i[9] vssa1 0.63fF
C636 user_analog_project_wrapper_empty_0/wbs_dat_o[8] vssa1 0.63fF
C637 user_analog_project_wrapper_empty_0/wbs_dat_i[8] vssa1 0.63fF
C638 user_analog_project_wrapper_empty_0/wbs_adr_i[8] vssa1 0.63fF
C639 user_analog_project_wrapper_empty_0/wbs_dat_o[7] vssa1 0.63fF
C640 user_analog_project_wrapper_empty_0/wbs_dat_i[7] vssa1 0.63fF
C641 user_analog_project_wrapper_empty_0/wbs_adr_i[7] vssa1 0.63fF
C642 user_analog_project_wrapper_empty_0/wbs_dat_o[6] vssa1 0.63fF
C643 user_analog_project_wrapper_empty_0/wbs_dat_i[6] vssa1 0.63fF
C644 user_analog_project_wrapper_empty_0/wbs_adr_i[6] vssa1 0.63fF
C645 user_analog_project_wrapper_empty_0/wbs_dat_o[5] vssa1 0.63fF
C646 user_analog_project_wrapper_empty_0/wbs_dat_i[5] vssa1 0.63fF
C647 user_analog_project_wrapper_empty_0/wbs_adr_i[5] vssa1 0.63fF
C648 user_analog_project_wrapper_empty_0/wbs_dat_o[4] vssa1 0.63fF
C649 user_analog_project_wrapper_empty_0/wbs_dat_i[4] vssa1 0.63fF
C650 user_analog_project_wrapper_empty_0/wbs_adr_i[4] vssa1 0.63fF
C651 user_analog_project_wrapper_empty_0/wbs_sel_i[3] vssa1 0.63fF
C652 user_analog_project_wrapper_empty_0/wbs_dat_o[3] vssa1 0.63fF
C653 user_analog_project_wrapper_empty_0/wbs_dat_i[3] vssa1 0.63fF
C654 user_analog_project_wrapper_empty_0/wbs_adr_i[3] vssa1 0.63fF
C655 user_analog_project_wrapper_empty_0/wbs_sel_i[2] vssa1 0.63fF
C656 user_analog_project_wrapper_empty_0/wbs_dat_o[2] vssa1 0.63fF
C657 user_analog_project_wrapper_empty_0/wbs_dat_i[2] vssa1 0.63fF
C658 user_analog_project_wrapper_empty_0/wbs_adr_i[2] vssa1 0.63fF
C659 user_analog_project_wrapper_empty_0/wbs_sel_i[1] vssa1 0.63fF
C660 user_analog_project_wrapper_empty_0/wbs_dat_o[1] vssa1 0.63fF
C661 user_analog_project_wrapper_empty_0/wbs_dat_i[1] vssa1 0.63fF
C662 user_analog_project_wrapper_empty_0/wbs_adr_i[1] vssa1 0.63fF
C663 user_analog_project_wrapper_empty_0/wbs_sel_i[0] vssa1 0.63fF
C664 user_analog_project_wrapper_empty_0/wbs_dat_o[0] vssa1 0.63fF
C665 user_analog_project_wrapper_empty_0/wbs_dat_i[0] vssa1 0.63fF
C666 user_analog_project_wrapper_empty_0/wbs_adr_i[0] vssa1 0.63fF
C667 user_analog_project_wrapper_empty_0/wbs_we_i vssa1 0.63fF
C668 user_analog_project_wrapper_empty_0/wbs_stb_i vssa1 0.63fF
C669 user_analog_project_wrapper_empty_0/wbs_cyc_i vssa1 0.63fF
C670 user_analog_project_wrapper_empty_0/wbs_ack_o vssa1 0.63fF
C671 user_analog_project_wrapper_empty_0/wb_rst_i vssa1 0.63fF
C672 user_analog_project_wrapper_empty_0/wb_clk_i vssa1 0.63fF
.ends

