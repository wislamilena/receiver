* SPICE3 file created from detV2.ext - technology: sky130A

.subckt detV2 din db do GND
X0 do bot_cin GND sky130_fd_pr__res_xhigh_po w=350000u l=1.86e+07u
X1 din bot_cin sky130_fd_pr__cap_mim_m3_1 l=8.7e+07u w=8.7e+07u
X2 do GND sky130_fd_pr__cap_mim_m3_1 l=8.7e+07u w=8.7e+07u
X3 GND db bot_cin GND sky130_fd_pr__nfet_01v8 w=2.25e+07u l=150000u
C0 bot_cin db 0.01fF
C1 bot_cin din 95.62fF
C2 din GND 5.43fF
C3 db GND 16.77fF
C4 do GND 126.12fF
C5 bot_cin GND 113.90fF **FLOATING
.ends
