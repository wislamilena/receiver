magic
tech sky130A
magscale 1 2
timestamp 1647304853
<< error_p >>
rect -11081 3200 -11021 9400
rect -11001 3200 -10941 9400
rect -4789 3200 -4729 9400
rect -4709 3200 -4649 9400
rect 1503 3200 1563 9400
rect 1583 3200 1643 9400
rect 7795 3200 7855 9400
rect 7875 3200 7935 9400
rect 14087 3200 14147 9400
rect 14167 3200 14227 9400
rect -11081 -3100 -11021 3100
rect -11001 -3100 -10941 3100
rect -4789 -3100 -4729 3100
rect -4709 -3100 -4649 3100
rect 1503 -3100 1563 3100
rect 1583 -3100 1643 3100
rect 7795 -3100 7855 3100
rect 7875 -3100 7935 3100
rect 14087 -3100 14147 3100
rect 14167 -3100 14227 3100
rect -11081 -9400 -11021 -3200
rect -11001 -9400 -10941 -3200
rect -4789 -9400 -4729 -3200
rect -4709 -9400 -4649 -3200
rect 1503 -9400 1563 -3200
rect 1583 -9400 1643 -3200
rect 7795 -9400 7855 -3200
rect 7875 -9400 7935 -3200
rect 14087 -9400 14147 -3200
rect 14167 -9400 14227 -3200
<< metal3 >>
rect -17293 9372 -11021 9400
rect -17293 3228 -11105 9372
rect -11041 3228 -11021 9372
rect -17293 3200 -11021 3228
rect -11001 9372 -4729 9400
rect -11001 3228 -4813 9372
rect -4749 3228 -4729 9372
rect -11001 3200 -4729 3228
rect -4709 9372 1563 9400
rect -4709 3228 1479 9372
rect 1543 3228 1563 9372
rect -4709 3200 1563 3228
rect 1583 9372 7855 9400
rect 1583 3228 7771 9372
rect 7835 3228 7855 9372
rect 1583 3200 7855 3228
rect 7875 9372 14147 9400
rect 7875 3228 14063 9372
rect 14127 3228 14147 9372
rect 7875 3200 14147 3228
rect 14167 9372 20439 9400
rect 14167 3228 20355 9372
rect 20419 3228 20439 9372
rect 14167 3200 20439 3228
rect -17293 3072 -11021 3100
rect -17293 -3072 -11105 3072
rect -11041 -3072 -11021 3072
rect -17293 -3100 -11021 -3072
rect -11001 3072 -4729 3100
rect -11001 -3072 -4813 3072
rect -4749 -3072 -4729 3072
rect -11001 -3100 -4729 -3072
rect -4709 3072 1563 3100
rect -4709 -3072 1479 3072
rect 1543 -3072 1563 3072
rect -4709 -3100 1563 -3072
rect 1583 3072 7855 3100
rect 1583 -3072 7771 3072
rect 7835 -3072 7855 3072
rect 1583 -3100 7855 -3072
rect 7875 3072 14147 3100
rect 7875 -3072 14063 3072
rect 14127 -3072 14147 3072
rect 7875 -3100 14147 -3072
rect 14167 3072 20439 3100
rect 14167 -3072 20355 3072
rect 20419 -3072 20439 3072
rect 14167 -3100 20439 -3072
rect -17293 -3228 -11021 -3200
rect -17293 -9372 -11105 -3228
rect -11041 -9372 -11021 -3228
rect -17293 -9400 -11021 -9372
rect -11001 -3228 -4729 -3200
rect -11001 -9372 -4813 -3228
rect -4749 -9372 -4729 -3228
rect -11001 -9400 -4729 -9372
rect -4709 -3228 1563 -3200
rect -4709 -9372 1479 -3228
rect 1543 -9372 1563 -3228
rect -4709 -9400 1563 -9372
rect 1583 -3228 7855 -3200
rect 1583 -9372 7771 -3228
rect 7835 -9372 7855 -3228
rect 1583 -9400 7855 -9372
rect 7875 -3228 14147 -3200
rect 7875 -9372 14063 -3228
rect 14127 -9372 14147 -3228
rect 7875 -9400 14147 -9372
rect 14167 -3228 20439 -3200
rect 14167 -9372 20355 -3228
rect 20419 -9372 20439 -3228
rect 14167 -9400 20439 -9372
<< via3 >>
rect -11105 3228 -11041 9372
rect -4813 3228 -4749 9372
rect 1479 3228 1543 9372
rect 7771 3228 7835 9372
rect 14063 3228 14127 9372
rect 20355 3228 20419 9372
rect -11105 -3072 -11041 3072
rect -4813 -3072 -4749 3072
rect 1479 -3072 1543 3072
rect 7771 -3072 7835 3072
rect 14063 -3072 14127 3072
rect 20355 -3072 20419 3072
rect -11105 -9372 -11041 -3228
rect -4813 -9372 -4749 -3228
rect 1479 -9372 1543 -3228
rect 7771 -9372 7835 -3228
rect 14063 -9372 14127 -3228
rect 20355 -9372 20419 -3228
<< mimcap >>
rect -17193 9260 -11193 9300
rect -17193 3340 -14785 9260
rect -13601 3340 -11193 9260
rect -17193 3300 -11193 3340
rect -10901 9260 -4901 9300
rect -10901 3340 -8493 9260
rect -7309 3340 -4901 9260
rect -10901 3300 -4901 3340
rect -4609 9260 1391 9300
rect -4609 3340 -2201 9260
rect -1017 3340 1391 9260
rect -4609 3300 1391 3340
rect 1683 9260 7683 9300
rect 1683 3340 4091 9260
rect 5275 3340 7683 9260
rect 1683 3300 7683 3340
rect 7975 9260 13975 9300
rect 7975 3340 10383 9260
rect 11567 3340 13975 9260
rect 7975 3300 13975 3340
rect 14267 9260 20267 9300
rect 14267 3340 16675 9260
rect 17859 3340 20267 9260
rect 14267 3300 20267 3340
rect -17193 2960 -11193 3000
rect -17193 -2960 -14785 2960
rect -13601 -2960 -11193 2960
rect -17193 -3000 -11193 -2960
rect -10901 2960 -4901 3000
rect -10901 -2960 -8493 2960
rect -7309 -2960 -4901 2960
rect -10901 -3000 -4901 -2960
rect -4609 2960 1391 3000
rect -4609 -2960 -2201 2960
rect -1017 -2960 1391 2960
rect -4609 -3000 1391 -2960
rect 1683 2960 7683 3000
rect 1683 -2960 4091 2960
rect 5275 -2960 7683 2960
rect 1683 -3000 7683 -2960
rect 7975 2960 13975 3000
rect 7975 -2960 10383 2960
rect 11567 -2960 13975 2960
rect 7975 -3000 13975 -2960
rect 14267 2960 20267 3000
rect 14267 -2960 16675 2960
rect 17859 -2960 20267 2960
rect 14267 -3000 20267 -2960
rect -17193 -3340 -11193 -3300
rect -17193 -9260 -14785 -3340
rect -13601 -9260 -11193 -3340
rect -17193 -9300 -11193 -9260
rect -10901 -3340 -4901 -3300
rect -10901 -9260 -8493 -3340
rect -7309 -9260 -4901 -3340
rect -10901 -9300 -4901 -9260
rect -4609 -3340 1391 -3300
rect -4609 -9260 -2201 -3340
rect -1017 -9260 1391 -3340
rect -4609 -9300 1391 -9260
rect 1683 -3340 7683 -3300
rect 1683 -9260 4091 -3340
rect 5275 -9260 7683 -3340
rect 1683 -9300 7683 -9260
rect 7975 -3340 13975 -3300
rect 7975 -9260 10383 -3340
rect 11567 -9260 13975 -3340
rect 7975 -9300 13975 -9260
rect 14267 -3340 20267 -3300
rect 14267 -9260 16675 -3340
rect 17859 -9260 20267 -3340
rect 14267 -9300 20267 -9260
<< mimcapcontact >>
rect -14785 3340 -13601 9260
rect -8493 3340 -7309 9260
rect -2201 3340 -1017 9260
rect 4091 3340 5275 9260
rect 10383 3340 11567 9260
rect 16675 3340 17859 9260
rect -14785 -2960 -13601 2960
rect -8493 -2960 -7309 2960
rect -2201 -2960 -1017 2960
rect 4091 -2960 5275 2960
rect 10383 -2960 11567 2960
rect 16675 -2960 17859 2960
rect -14785 -9260 -13601 -3340
rect -8493 -9260 -7309 -3340
rect -2201 -9260 -1017 -3340
rect 4091 -9260 5275 -3340
rect 10383 -9260 11567 -3340
rect 16675 -9260 17859 -3340
<< metal4 >>
rect -11121 9372 -11025 9388
rect -14786 9260 -13600 9261
rect -14786 3340 -14785 9260
rect -13601 3340 -13600 9260
rect -14786 3339 -13600 3340
rect -11121 3228 -11105 9372
rect -11041 3228 -11025 9372
rect -4829 9372 -4733 9388
rect -8494 9260 -7308 9261
rect -8494 3340 -8493 9260
rect -7309 3340 -7308 9260
rect -8494 3339 -7308 3340
rect -11121 3212 -11025 3228
rect -4829 3228 -4813 9372
rect -4749 3228 -4733 9372
rect 1463 9372 1559 9388
rect -2202 9260 -1016 9261
rect -2202 3340 -2201 9260
rect -1017 3340 -1016 9260
rect -2202 3339 -1016 3340
rect -4829 3212 -4733 3228
rect 1463 3228 1479 9372
rect 1543 3228 1559 9372
rect 7755 9372 7851 9388
rect 4090 9260 5276 9261
rect 4090 3340 4091 9260
rect 5275 3340 5276 9260
rect 4090 3339 5276 3340
rect 1463 3212 1559 3228
rect 7755 3228 7771 9372
rect 7835 3228 7851 9372
rect 14047 9372 14143 9388
rect 10382 9260 11568 9261
rect 10382 3340 10383 9260
rect 11567 3340 11568 9260
rect 10382 3339 11568 3340
rect 7755 3212 7851 3228
rect 14047 3228 14063 9372
rect 14127 3228 14143 9372
rect 20339 9372 20435 9388
rect 16674 9260 17860 9261
rect 16674 3340 16675 9260
rect 17859 3340 17860 9260
rect 16674 3339 17860 3340
rect 14047 3212 14143 3228
rect 20339 3228 20355 9372
rect 20419 3228 20435 9372
rect 20339 3212 20435 3228
rect -11121 3072 -11025 3088
rect -14786 2960 -13600 2961
rect -14786 -2960 -14785 2960
rect -13601 -2960 -13600 2960
rect -14786 -2961 -13600 -2960
rect -11121 -3072 -11105 3072
rect -11041 -3072 -11025 3072
rect -4829 3072 -4733 3088
rect -8494 2960 -7308 2961
rect -8494 -2960 -8493 2960
rect -7309 -2960 -7308 2960
rect -8494 -2961 -7308 -2960
rect -11121 -3088 -11025 -3072
rect -4829 -3072 -4813 3072
rect -4749 -3072 -4733 3072
rect 1463 3072 1559 3088
rect -2202 2960 -1016 2961
rect -2202 -2960 -2201 2960
rect -1017 -2960 -1016 2960
rect -2202 -2961 -1016 -2960
rect -4829 -3088 -4733 -3072
rect 1463 -3072 1479 3072
rect 1543 -3072 1559 3072
rect 7755 3072 7851 3088
rect 4090 2960 5276 2961
rect 4090 -2960 4091 2960
rect 5275 -2960 5276 2960
rect 4090 -2961 5276 -2960
rect 1463 -3088 1559 -3072
rect 7755 -3072 7771 3072
rect 7835 -3072 7851 3072
rect 14047 3072 14143 3088
rect 10382 2960 11568 2961
rect 10382 -2960 10383 2960
rect 11567 -2960 11568 2960
rect 10382 -2961 11568 -2960
rect 7755 -3088 7851 -3072
rect 14047 -3072 14063 3072
rect 14127 -3072 14143 3072
rect 20339 3072 20435 3088
rect 16674 2960 17860 2961
rect 16674 -2960 16675 2960
rect 17859 -2960 17860 2960
rect 16674 -2961 17860 -2960
rect 14047 -3088 14143 -3072
rect 20339 -3072 20355 3072
rect 20419 -3072 20435 3072
rect 20339 -3088 20435 -3072
rect -11121 -3228 -11025 -3212
rect -14786 -3340 -13600 -3339
rect -14786 -9260 -14785 -3340
rect -13601 -9260 -13600 -3340
rect -14786 -9261 -13600 -9260
rect -11121 -9372 -11105 -3228
rect -11041 -9372 -11025 -3228
rect -4829 -3228 -4733 -3212
rect -8494 -3340 -7308 -3339
rect -8494 -9260 -8493 -3340
rect -7309 -9260 -7308 -3340
rect -8494 -9261 -7308 -9260
rect -11121 -9388 -11025 -9372
rect -4829 -9372 -4813 -3228
rect -4749 -9372 -4733 -3228
rect 1463 -3228 1559 -3212
rect -2202 -3340 -1016 -3339
rect -2202 -9260 -2201 -3340
rect -1017 -9260 -1016 -3340
rect -2202 -9261 -1016 -9260
rect -4829 -9388 -4733 -9372
rect 1463 -9372 1479 -3228
rect 1543 -9372 1559 -3228
rect 7755 -3228 7851 -3212
rect 4090 -3340 5276 -3339
rect 4090 -9260 4091 -3340
rect 5275 -9260 5276 -3340
rect 4090 -9261 5276 -9260
rect 1463 -9388 1559 -9372
rect 7755 -9372 7771 -3228
rect 7835 -9372 7851 -3228
rect 14047 -3228 14143 -3212
rect 10382 -3340 11568 -3339
rect 10382 -9260 10383 -3340
rect 11567 -9260 11568 -3340
rect 10382 -9261 11568 -9260
rect 7755 -9388 7851 -9372
rect 14047 -9372 14063 -3228
rect 14127 -9372 14143 -3228
rect 20339 -3228 20435 -3212
rect 16674 -3340 17860 -3339
rect 16674 -9260 16675 -3340
rect 17859 -9260 17860 -3340
rect 16674 -9261 17860 -9260
rect 14047 -9388 14143 -9372
rect 20339 -9372 20355 -3228
rect 20419 -9372 20435 -3228
rect 20339 -9388 20435 -9372
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 14167 3200 20367 9400
string parameters w 30.0 l 30.0 val 920.4 carea 1.00 cperi 0.17 nx 5.5 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 20
string library sky130
<< end >>
