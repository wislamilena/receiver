magic
tech sky130A
magscale 1 2
timestamp 1647304558
<< error_p >>
rect -29 2322 29 2328
rect -29 2288 -17 2322
rect -29 2282 29 2288
rect -29 -2288 29 -2282
rect -29 -2322 -17 -2288
rect -29 -2328 29 -2322
<< nmos >>
rect -15 -2250 15 2250
<< ndiff >>
rect -73 2238 -15 2250
rect -73 -2238 -61 2238
rect -27 -2238 -15 2238
rect -73 -2250 -15 -2238
rect 15 2238 73 2250
rect 15 -2238 27 2238
rect 61 -2238 73 2238
rect 15 -2250 73 -2238
<< ndiffc >>
rect -61 -2238 -27 2238
rect 27 -2238 61 2238
<< poly >>
rect -33 2322 33 2338
rect -33 2288 -17 2322
rect 17 2288 33 2322
rect -33 2272 33 2288
rect -15 2250 15 2272
rect -15 -2272 15 -2250
rect -33 -2288 33 -2272
rect -33 -2322 -17 -2288
rect 17 -2322 33 -2288
rect -33 -2338 33 -2322
<< polycont >>
rect -17 2288 17 2322
rect -17 -2322 17 -2288
<< locali >>
rect -33 2288 -17 2322
rect 17 2288 33 2322
rect -61 2238 -27 2254
rect -61 -2254 -27 -2238
rect 27 2238 61 2254
rect 27 -2254 61 -2238
rect -33 -2322 -17 -2288
rect 17 -2322 33 -2288
<< viali >>
rect -17 2288 17 2322
rect -61 -2238 -27 2238
rect 27 -2238 61 2238
rect -17 -2322 17 -2288
<< metal1 >>
rect -29 2322 29 2328
rect -29 2288 -17 2322
rect 17 2288 29 2322
rect -29 2282 29 2288
rect -67 2238 -21 2250
rect -67 -2238 -61 2238
rect -27 -2238 -21 2238
rect -67 -2250 -21 -2238
rect 21 2238 67 2250
rect 21 -2238 27 2238
rect 61 -2238 67 2238
rect 21 -2250 67 -2238
rect -29 -2288 29 -2282
rect -29 -2322 -17 -2288
rect 17 -2322 29 -2288
rect -29 -2328 29 -2322
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 22.5 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 1 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
