*************************************************************************************
.TITLE TEST BENCH DETECTOR

.LIB /edatools/pdks/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt
.INCLUDE /home/wisla/sky130_skel/Myschematics/Receptor/askMod.spice
.INCLUDE /home/wisla/sky130_skel/Myschematics/Receptor/my_chip/caravel_user_project_analog/xschem/detector.spice

* CALL SUBCIRCUIT
Xdet din db do GND detectorPassivo
Xask din GND askMod
Vb db GND 1

.TRAN 1p 250n
.GLOBAL GND
.END
