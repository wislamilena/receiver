* SPICE3 file created from otaV5.ext - technology: sky130A

.subckt otaV5 Inp Inn Vout Ib cltop Vp Vn
X0 Vn a_6890_1010# a_6890_750# Vn sky130_fd_pr__nfet_01v8 w=800000u l=4e+06u
X1 a_7570_1796# Inp a_6890_1010# Vp sky130_fd_pr__pfet_01v8 w=1.7e+06u l=2e+06u
X2 Vn a_8070_1014# a_8070_1014# Vn sky130_fd_pr__nfet_01v8 w=800000u l=4e+06u
X3 Vn a_6890_1010# a_6890_1010# Vn sky130_fd_pr__nfet_01v8 w=800000u l=4e+06u
X4 Vp a_6890_750# Vout Vp sky130_fd_pr__pfet_01v8 w=1.4e+06u l=1e+06u
X5 Vp Ib a_7570_1796# Vp sky130_fd_pr__pfet_01v8 w=5e+06u l=4e+06u
X6 cltop Vout sky130_fd_pr__cap_mim_m3_1 l=3.2e+07u w=3.2e+07u
X7 Vn a_8070_1014# Vout Vn sky130_fd_pr__nfet_01v8 w=800000u l=4e+06u
X8 Vp a_6890_750# a_6890_750# Vp sky130_fd_pr__pfet_01v8 w=1.4e+06u l=1e+06u
X9 a_8070_1014# Inn a_7570_1796# Vp sky130_fd_pr__pfet_01v8 w=1.7e+06u l=2e+06u
X10 Vp Ib Ib Vp sky130_fd_pr__pfet_01v8 w=5e+06u l=4e+06u
C0 a_6890_1010# a_6890_750# 0.44fF
C1 Inn a_8070_1014# 0.03fF
C2 Inn Inp 0.37fF
C3 a_8070_1014# a_6890_750# 0.07fF
C4 Inp Vp 0.17fF
C5 a_8070_1014# Vout 0.09fF
C6 Inp Ib 0.08fF
C7 a_6890_750# Vp 0.09fF
C8 cltop Vout 15.77fF
C9 a_8070_1014# a_6890_1010# 0.01fF
C10 Inp a_6890_1010# 0.16fF
C11 Inn Ib 0.11fF
C12 a_7570_1796# Vp 0.01fF
C13 Ib Vp 0.27fF
C14 Vout Vp 0.03fF
C15 Inn a_6890_1010# 0.22fF
C16 a_6890_750# Vout 1.07fF
C17 cltop Vn 1.16fF
C18 Vout Vn 28.38fF
C19 Inn Vn 2.75fF
C20 Inp Vn 7.19fF
C21 Ib Vn 7.73fF
C22 Vp Vn 31.12fF
C23 a_8070_1014# Vn 2.45fF **FLOATING
C24 a_6890_1010# Vn 2.61fF **FLOATING
C25 a_6890_750# Vn 2.36fF **FLOATING
C26 a_7570_1796# Vn 0.10fF **FLOATING
.ends
