** sch_path: /home/wisla/sky130_skel/Myschematics/Receptor/EnvelopeDetector/tb_detectorASK.sch
**.subckt tb_detectorASK
X1 ask vb GND out detectorPassivo
V1 vb GND 0.9
X2 ask GND askMod
**** begin user architecture code


.tran 1e-10 100u
.control
 run
 plot out
.endc



.lib /edatools/pdks/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/sky130.lib.spice tt

**** end user architecture code
**.ends

* expanding   symbol:  /home/wisla/sky130_skel/Myschematics/detectorPassivo.sym # of pins=4
** sym_path: /home/wisla/sky130_skel/Myschematics/detectorPassivo.sym
** sch_path: /home/wisla/sky130_skel/Myschematics/detectorPassivo.sch
.subckt detectorPassivo  din dB ground do
*.ipin din
*.ipin dB
*.opin do
*.iopin gnd
XM1 net1 dB gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC3 do gnd sky130_fd_pr__cap_mim_m3_2 W=22 L=22 VM=1 m=1
XR2 do net1 gnd sky130_fd_pr__res_xhigh_po W=0.35 L=17.5 mult=1 m=1
XC1 din net1 sky130_fd_pr__cap_mim_m3_2 W=87 L=87 VM=1 m=1
.ends


* expanding   symbol:  /home/wisla/sky130_skel/Myschematics/Receptor/EnvelopeDetector/askMod.sym #
*+ of pins=2
** sym_path: /home/wisla/sky130_skel/Myschematics/Receptor/EnvelopeDetector/askMod.sym
** sch_path: /home/wisla/sky130_skel/Myschematics/Receptor/EnvelopeDetector/askMod.sch
.subckt askMod  ask ground
*.opin ask
*.iopin gnd
XM2 carrier DS ask gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
R1 ask gnd 10 m=1
V3 DS gnd PULSE(0 1.8 100n 100n 100n 32u 64u)
V1 carrier gnd sin(0 500m 2e9)
.ends

.GLOBAL GND
.end
