* NGSPICE file created from otaV5.ext - technology: sky130A

.subckt otaV5 Inp Inn Vout Ib cltop Vp Vn
X0 Vn.t3 a_6890_1010.t3 a_6890_750.t2 Vn sky130_fd_pr__nfet_01v8 w=800000u l=4e+06u
X1 a_7570_1796.t2 Inp.t0 a_6890_1010.t0 Vp.t6 sky130_fd_pr__pfet_01v8 w=1.7e+06u l=2e+06u
X2 Vn.t0 a_8070_1014.t1 a_8070_1014.t2 Vn sky130_fd_pr__nfet_01v8 w=800000u l=4e+06u
X3 Vn.t2 a_6890_1010.t1 a_6890_1010.t2 Vn sky130_fd_pr__nfet_01v8 w=800000u l=4e+06u
X4 Vp.t5 a_6890_750.t3 Vout.t0 Vp.t3 sky130_fd_pr__pfet_01v8 w=1.4e+06u l=1e+06u
X5 Vp.t2 Ib.t0 a_7570_1796.t1 Vp.t1 sky130_fd_pr__pfet_01v8 w=5e+06u l=4e+06u
X6 cltop.t0 Vout.t1 sky130_fd_pr__cap_mim_m3_1 l=3.2e+07u w=3.2e+07u
X7 Vn.t1 a_8070_1014.t3 Vout.t2 Vn sky130_fd_pr__nfet_01v8 w=800000u l=4e+06u
X8 Vp.t4 a_6890_750.t0 a_6890_750.t1 Vp.t3 sky130_fd_pr__pfet_01v8 w=1.4e+06u l=1e+06u
X9 a_8070_1014.t0 Inn.t0 a_7570_1796.t0 Vp.t0 sky130_fd_pr__pfet_01v8 w=1.7e+06u l=2e+06u
X10 Vp Ib Ib Vp sky130_fd_pr__pfet_01v8 w=5e+06u l=4e+06u
R0 a_6890_1010.t0 a_6890_1010.n0 195.921
R1 a_6890_1010.n0 a_6890_1010.t1 92.645
R2 a_6890_1010.n0 a_6890_1010.t2 69.562
R3 a_6890_1010.t1 a_6890_1010.t3 10.845
R4 a_6890_750.n0 a_6890_750.t0 207.335
R5 a_6890_750.t0 a_6890_750.t3 91.58
R6 a_6890_750.n0 a_6890_750.t2 80.953
R7 a_6890_750.t1 a_6890_750.n0 63.038
R8 Vn.n1 Vn.t2 84.412
R9 Vn.n2 Vn.n0 65.938
R10 Vn.n0 Vn.t0 65.166
R11 Vn.n2 Vn.n1 63.208
R12 Vn.n0 Vn.t1 38.25
R13 Vn.n1 Vn.t3 38.25
R14 Vn Vn.n2 0.006
R15 Inp Inp.t0 27.195
R16 a_7570_1796.t1 a_7570_1796.n0 873.24
R17 a_7570_1796.n0 a_7570_1796.t0 29.55
R18 a_7570_1796.n0 a_7570_1796.t2 28.391
R19 Vp.n1 Vp.t2 1996.51
R20 Vp.n2 Vp.n1 722.838
R21 Vp.n2 Vp.t4 598.495
R22 Vp.t4 Vp.t5 434.506
R23 Vp.n0 Vp.t1 322.249
R24 Vp.n0 Vp.t3 306.762
R25 Vp.t0 Vp.t6 297.827
R26 Vp.t1 Vp.t0 119.131
R27 Vp.n1 Vp.n0 3.566
R28 Vp Vp.n2 0.145
R29 a_8070_1014.t0 a_8070_1014.n0 304.285
R30 a_8070_1014.n0 a_8070_1014.t1 85.41
R31 a_8070_1014.n0 a_8070_1014.t2 59.814
R32 a_8070_1014.t1 a_8070_1014.t3 10.845
R33 Vout.n0 Vout.t0 210.109
R34 Vout.n0 Vout.t1 166.261
R35 Vout.n1 Vout.t2 56.397
R36 Vout Vout.n1 0.067
R37 Vout.n1 Vout.n0 0.001
R38 Ib Ib.n1 840.712
R39 Ib Ib.n0 84.078
R40 Ib.n0 Ib.t0 68.685
R41 cltop cltop.t0 0.054
R42 Inn.n0 Inn.t0 20.485
R43 Inn.n0 Inn 4.357
R44 Inn Inn.n0 2.614
C0 Vp Ib 0.27fF
C1 Inp Inn 0.37fF
C2 Ib Inn 0.11fF
C3 Vp Vout 0.03fF
C4 Inp Vp 0.17fF
C5 cltop Vout 15.92fF
C6 Inp Ib 0.08fF
.ends

