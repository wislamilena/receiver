magic
tech sky130A
magscale 1 2
timestamp 1654529013
<< nmos >>
rect 2246 1280 2276 3080
<< ndiff >>
rect 2170 2963 2246 3080
rect 2170 2911 2180 2963
rect 2214 2911 2246 2963
rect 2170 2763 2246 2911
rect 2170 2711 2180 2763
rect 2214 2711 2246 2763
rect 2170 2563 2246 2711
rect 2170 2511 2180 2563
rect 2214 2511 2246 2563
rect 2170 2363 2246 2511
rect 2170 2311 2180 2363
rect 2214 2311 2246 2363
rect 2170 2163 2246 2311
rect 2170 2111 2180 2163
rect 2214 2111 2246 2163
rect 2170 1963 2246 2111
rect 2170 1911 2180 1963
rect 2214 1911 2246 1963
rect 2170 1763 2246 1911
rect 2170 1711 2180 1763
rect 2214 1711 2246 1763
rect 2170 1563 2246 1711
rect 2170 1511 2180 1563
rect 2214 1511 2246 1563
rect 2170 1362 2246 1511
rect 2170 1310 2180 1362
rect 2214 1310 2246 1362
rect 2170 1280 2246 1310
rect 2276 2962 2352 3080
rect 2276 2910 2310 2962
rect 2344 2910 2352 2962
rect 2276 2762 2352 2910
rect 2276 2710 2310 2762
rect 2344 2710 2352 2762
rect 2276 2562 2352 2710
rect 2276 2510 2310 2562
rect 2344 2510 2352 2562
rect 2276 2362 2352 2510
rect 2276 2310 2310 2362
rect 2344 2310 2352 2362
rect 2276 2162 2352 2310
rect 2276 2110 2310 2162
rect 2344 2110 2352 2162
rect 2276 1962 2352 2110
rect 2276 1910 2310 1962
rect 2344 1910 2352 1962
rect 2276 1762 2352 1910
rect 2276 1710 2310 1762
rect 2344 1710 2352 1762
rect 2276 1562 2352 1710
rect 2276 1510 2310 1562
rect 2344 1510 2352 1562
rect 2276 1362 2352 1510
rect 2276 1310 2310 1362
rect 2344 1310 2352 1362
rect 2276 1280 2352 1310
<< ndiffc >>
rect 2180 2911 2214 2963
rect 2180 2711 2214 2763
rect 2180 2511 2214 2563
rect 2180 2311 2214 2363
rect 2180 2111 2214 2163
rect 2180 1911 2214 1963
rect 2180 1711 2214 1763
rect 2180 1511 2214 1563
rect 2180 1310 2214 1362
rect 2310 2910 2344 2962
rect 2310 2710 2344 2762
rect 2310 2510 2344 2562
rect 2310 2310 2344 2362
rect 2310 2110 2344 2162
rect 2310 1910 2344 1962
rect 2310 1710 2344 1762
rect 2310 1510 2344 1562
rect 2310 1310 2344 1362
<< psubdiff >>
rect 2352 3042 2428 3080
rect 2352 2990 2364 3042
rect 2398 2990 2428 3042
rect 2352 2842 2428 2990
rect 2352 2790 2364 2842
rect 2398 2790 2428 2842
rect 2352 2642 2428 2790
rect 2352 2590 2364 2642
rect 2398 2590 2428 2642
rect 2352 2442 2428 2590
rect 2352 2390 2364 2442
rect 2398 2390 2428 2442
rect 2352 2242 2428 2390
rect 2352 2190 2364 2242
rect 2398 2190 2428 2242
rect 2352 2042 2428 2190
rect 2352 1990 2364 2042
rect 2398 1990 2428 2042
rect 2352 1842 2428 1990
rect 2352 1790 2364 1842
rect 2398 1790 2428 1842
rect 2352 1642 2428 1790
rect 2352 1590 2364 1642
rect 2398 1590 2428 1642
rect 2352 1442 2428 1590
rect 2352 1390 2364 1442
rect 2398 1390 2428 1442
rect 2352 1280 2428 1390
<< psubdiffcont >>
rect 2364 2990 2398 3042
rect 2364 2790 2398 2842
rect 2364 2590 2398 2642
rect 2364 2390 2398 2442
rect 2364 2190 2398 2242
rect 2364 1990 2398 2042
rect 2364 1790 2398 1842
rect 2364 1590 2398 1642
rect 2364 1390 2398 1442
<< poly >>
rect 2246 3080 2276 3130
rect 2246 1236 2276 1280
rect 2246 1200 2432 1236
rect 2246 1034 2278 1200
rect 2398 1034 2432 1200
rect 2246 1000 2432 1034
<< polycont >>
rect 2278 1034 2398 1200
<< xpolycontact >>
rect 2690 3898 2760 4426
rect 2690 -130 2760 398
<< xpolyres >>
rect 2690 398 2760 3898
<< locali >>
rect 2170 4116 2690 4166
rect 2170 3060 2218 4116
rect 2300 3410 2414 3418
rect 2300 3316 2314 3410
rect 2400 3316 2414 3410
rect 2300 3310 2414 3316
rect 2332 3060 2380 3310
rect 2170 2963 2220 3060
rect 2170 2911 2180 2963
rect 2214 2911 2220 2963
rect 2170 2763 2220 2911
rect 2170 2711 2180 2763
rect 2214 2711 2220 2763
rect 2170 2563 2220 2711
rect 2170 2511 2180 2563
rect 2214 2511 2220 2563
rect 2170 2370 2220 2511
rect 2040 2363 2220 2370
rect 2040 2330 2180 2363
rect 2040 2240 2060 2330
rect 2130 2311 2180 2330
rect 2214 2311 2220 2363
rect 2130 2240 2220 2311
rect 2040 2163 2220 2240
rect 2040 2111 2180 2163
rect 2214 2111 2220 2163
rect 2040 2030 2220 2111
rect 2040 1940 2060 2030
rect 2130 1963 2220 2030
rect 2130 1940 2180 1963
rect 2040 1911 2180 1940
rect 2214 1911 2220 1963
rect 2040 1910 2220 1911
rect 2170 1763 2220 1910
rect 2170 1711 2180 1763
rect 2214 1711 2220 1763
rect 2170 1563 2220 1711
rect 2170 1511 2180 1563
rect 2214 1511 2220 1563
rect 2170 1362 2220 1511
rect 2170 1310 2180 1362
rect 2214 1310 2220 1362
rect 2170 1290 2220 1310
rect 2300 3042 2410 3060
rect 2300 2990 2364 3042
rect 2398 2990 2410 3042
rect 2300 2962 2410 2990
rect 2300 2910 2310 2962
rect 2344 2910 2410 2962
rect 2300 2842 2410 2910
rect 2300 2790 2364 2842
rect 2398 2790 2410 2842
rect 2300 2762 2410 2790
rect 2300 2710 2310 2762
rect 2344 2710 2410 2762
rect 2300 2642 2410 2710
rect 2300 2590 2364 2642
rect 2398 2590 2410 2642
rect 2300 2562 2410 2590
rect 2300 2510 2310 2562
rect 2344 2510 2410 2562
rect 2300 2442 2410 2510
rect 2300 2390 2364 2442
rect 2398 2390 2410 2442
rect 2300 2362 2410 2390
rect 2300 2310 2310 2362
rect 2344 2310 2410 2362
rect 2300 2242 2410 2310
rect 2300 2190 2364 2242
rect 2398 2190 2410 2242
rect 2300 2162 2410 2190
rect 2300 2110 2310 2162
rect 2344 2110 2410 2162
rect 2300 2042 2410 2110
rect 2300 1990 2364 2042
rect 2398 1990 2410 2042
rect 2300 1962 2410 1990
rect 2300 1910 2310 1962
rect 2344 1910 2410 1962
rect 2300 1842 2410 1910
rect 2300 1790 2364 1842
rect 2398 1790 2410 1842
rect 2300 1762 2410 1790
rect 2300 1710 2310 1762
rect 2344 1710 2410 1762
rect 2300 1642 2410 1710
rect 2300 1590 2364 1642
rect 2398 1590 2410 1642
rect 2300 1562 2410 1590
rect 2300 1510 2310 1562
rect 2344 1510 2410 1562
rect 2300 1442 2410 1510
rect 2300 1390 2364 1442
rect 2398 1390 2410 1442
rect 2300 1362 2410 1390
rect 2300 1310 2310 1362
rect 2344 1310 2410 1362
rect 2300 1290 2410 1310
rect 2246 1200 2432 1236
rect 2246 1034 2278 1200
rect 2398 1034 2432 1200
rect 2246 1000 2432 1034
rect 2842 276 3210 358
rect 2842 232 2914 276
rect 2760 -34 2914 232
rect 2842 -46 2914 -34
rect 3150 -46 3210 276
rect 2842 -100 3210 -46
<< viali >>
rect 2314 3316 2400 3410
rect 2060 2240 2130 2330
rect 2060 1940 2130 2030
rect 2278 1034 2398 1200
rect 2914 -46 3150 276
<< metal1 >>
rect 2300 3410 2414 3418
rect 2300 3316 2314 3410
rect 2400 3316 2414 3410
rect 2300 3310 2414 3316
rect 2040 2330 2150 2370
rect 2040 2240 2060 2330
rect 2130 2240 2150 2330
rect 2040 2030 2150 2240
rect 2040 1940 2060 2030
rect 2130 1940 2150 2030
rect 2040 1910 2150 1940
rect 2246 1200 2432 1236
rect 2246 1034 2278 1200
rect 2398 1034 2432 1200
rect 2246 1000 2432 1034
rect 2842 276 3210 358
rect 2842 -46 2914 276
rect 3150 -46 3210 276
rect 2842 -100 3210 -46
<< via1 >>
rect 2314 3316 2400 3410
rect 2060 2240 2130 2330
rect 2060 1940 2130 2030
rect 2278 1034 2398 1200
rect 2914 -46 3150 276
<< metal2 >>
rect 2300 3410 2414 3418
rect 2300 3316 2314 3410
rect 2400 3316 2414 3410
rect 2300 3310 2414 3316
rect 2040 2330 2150 2370
rect 2040 2240 2060 2330
rect 2130 2240 2150 2330
rect 2040 2030 2150 2240
rect 2040 1940 2060 2030
rect 2130 1940 2150 2030
rect 2040 1910 2150 1940
rect 2246 1200 2432 1236
rect 2246 1034 2278 1200
rect 2398 1034 2432 1200
rect 2246 1000 2432 1034
rect 2842 276 3210 358
rect 2842 -46 2914 276
rect 3150 -46 3210 276
rect 2842 -100 3210 -46
<< via2 >>
rect 2314 3316 2400 3410
rect 2060 2240 2130 2330
rect 2060 1940 2130 2030
rect 2278 1034 2398 1200
rect 2914 -46 3150 276
<< metal3 >>
rect 8100 4966 8400 5002
rect 8100 4900 8132 4966
rect 2332 4800 8132 4900
rect 2332 3418 2394 4800
rect 8100 4748 8132 4800
rect 8368 4748 8400 4966
rect 8100 4698 8400 4748
rect 2300 3410 2414 3418
rect 2300 3316 2314 3410
rect 2400 3316 2414 3410
rect 2300 3310 2414 3316
rect 2040 2330 2150 2370
rect 2040 2240 2060 2330
rect 2130 2240 2150 2330
rect 2040 2030 2150 2240
rect 2040 1940 2060 2030
rect 2130 1940 2150 2030
rect 2040 1910 2150 1940
rect 2246 1200 2432 1236
rect 2246 1034 2278 1200
rect 2398 1034 2432 1200
rect 2246 1000 2432 1034
rect 2842 276 3210 358
rect 2842 -46 2914 276
rect 3150 -46 3210 276
rect 2842 -100 3210 -46
<< via3 >>
rect 8132 4748 8368 4966
rect 2060 2240 2130 2330
rect 2060 1940 2130 2030
rect 2278 1034 2398 1200
rect 2914 -46 3150 276
<< metal4 >>
rect -18058 2370 2024 14998
rect 8100 4966 8400 5002
rect 8100 4748 8132 4966
rect 8368 4748 8400 4966
rect 8100 4500 8400 4748
rect -18058 2330 2150 2370
rect -18058 2240 2060 2330
rect 2130 2240 2150 2330
rect -18058 2030 2150 2240
rect -18058 1940 2060 2030
rect 2130 1940 2150 2030
rect -18058 1910 2150 1940
rect -18058 -4976 2024 1910
rect 2246 1200 2432 1236
rect 2246 1034 2278 1200
rect 2398 1034 2432 1200
rect 2246 1000 2432 1034
rect 2300 -602 2372 1000
rect 2842 276 3210 358
rect 2842 -46 2914 276
rect 3150 -46 3210 276
rect 2842 -100 3210 -46
rect 3446 -360 8438 4500
rect 8328 -602 8518 -514
rect 2300 -672 8518 -602
rect 8328 -780 8518 -672
<< via4 >>
rect 2914 -46 3150 276
<< mimcap2 >>
rect -17002 6054 398 13372
rect -17002 2980 -15008 6054
rect -11984 2980 398 6054
rect -17002 -4028 398 2980
rect 3710 308 8110 4250
rect 3710 -60 3800 308
rect 5650 -60 8110 308
rect 3710 -150 8110 -60
<< mimcap2contact >>
rect -15008 2980 -11984 6054
rect 3800 -60 5650 308
<< metal5 >>
rect -20000 6054 -10006 6998
rect -20000 2980 -15008 6054
rect -11984 2980 -10006 6054
rect -20000 1998 -10006 2980
rect 5722 400 8440 402
rect 3268 358 8440 400
rect 2842 308 8440 358
rect 2842 276 3800 308
rect 2842 -46 2914 276
rect 3150 -46 3800 276
rect 2842 -60 3800 -46
rect 5650 -60 8440 308
rect 2842 -100 8440 -60
rect 3268 -152 8440 -100
<< labels >>
flabel metal5 -19580 2548 -18152 6054 0 FreeSans 4800 0 0 0 din
port 1 nsew
flabel locali 2300 2408 2338 2482 0 FreeSans 160 0 0 0 nbs
flabel metal5 2930 -50 3158 280 0 FreeSans 320 0 0 0 rc
flabel metal5 8126 -84 8378 246 0 FreeSans 1600 0 0 0 do
port 3 nsew
flabel metal4 8330 -780 8516 -516 0 FreeSans 480 0 0 0 db
port 2 nsew
flabel locali 2046 2096 2162 2194 0 FreeSans 160 0 0 0 nd
flabel metal4 8116 4748 8370 4972 0 FreeSans 480 0 0 0 GND
port 4 nsew
<< end >>
